��/  ���a��|[�{-r�#nl[m�v�{5��7MZ�|b��}�"�8LX��(�Z�ʱO�'�Z�i�%��7�B�^��8$�0������P�5#�E��w�9�@�\V1����,��r\��>!���N,��
po�I�;ط�&[��� �AuxN�����h4�*�> ��c>%$;��]�q��3p����.���\06D橧��@hH�U��QJ6eN��f�2;Al�͓�Ƥ�p�-�}Д�)U��U!����\tØ��}sz�.����2�ȴ�l H��8~�u�V��S���QA.��-Rӊ"�d7�_U���5�N�!_�����T��$��c(iX��(d����i�`i #���0�'> %lz�},/�P��/�dy�ԲU��o����P��/���1DA,��,	�d���'������|��-;Mퟻ$��vU���O�e��M����3�7T�ir�V��
�˫Tn3��H���ϢƖC1���*LHk��}E���V�а5;%
�o�Ps&2�O��Q����שv�E^tJ�sg耼A�20y0��h�3��K9���R.��^����MᾸ={"��Xc�r�e�Ǹ��ߢ[z�U�s}"�H���+��H��ې`ѱ.��XP�)�4���cqs�����x�����O�Ҕ0V� ��ըH#=�~���E_֌��/�>l�Y�[L-�;��	���.)"p�J-����+ѷ�6X�H@��E1rF���)/�C�o~8MmL�-�'�:�hG9�:Y��(ma�[�?�w���Co&��*���>w��c6p���v[�}������8�����址�PBW,㎺VCv*b�<3N�)=���.ŗ*Ɛ��P©͔��Kd��=��:���'ʮ�펧U�'���u�p+��a�u�7�~�a̿��daDRUs��]P��y�b��b$erF�� ;�l(H\�3���"�5`aA��#�"FYf�N��z�4���3iW��O-K��Q�*8�9߰X[�o@p��d^�U�h���!rJ��Ѭ�Gø�/`ݏh5���Wz�N�z��bP�?>�,�I��O��M�(BvP�A`�I������>?�J���X&oO�o��������Aq����s[OJ��M��Oj�}1�%֤��)��RI��p���!�K�c��)^��mn]JՋ��q��/|/#rT�t㯍�u��ҧ%�j�N�͹�0&�/�5j#1z�v�͇�ŋ ٿ��f�rO>�|����k����Q�2L�rb�4�x�6��/Sh�� ��#���I��'�n�tYޱ=l�^l�]sR�����<�x�����Y���q�� =O���-��gH��)	(���Ϭ�jS-�++���;�+�B�O�%�d^B����=ot|��׏o��ڎ���N������k�7�]o��E7:�9h�埈b�B�N���`<��,�$N�+؈�7�?�7Qo��.���ֹѸ¾��s[03ԛ���h��1�P6fD1ab����V?&���j�7-d�v��gm��E1���,]��r�5{�@H����d�����1톡R��V��t��=!����i-�}W�T� A��߷���6���s�q�0������c�`������+ ����Y�\�P�m�Z�c��e97~@����3����7�A��4�D���dq¶q��w����LM��&�G����O�<���}�Mv���_��XQi��27�e�����;��Mkr�#9�7a��N;�H �4'��+�e�&$W�{��HKCX�_���UC��g@���+b��zH�Y�" �l������Y�ޠ��[�r,pZH�O���߮��-FW���6����f�>:�eCP�y��6	EC�Z[�u��=���[cz��+��ߛ.�K�@�D2s;D���E��"oM�t��R�j��UJ�[o$�h]�X,���{HqrR��b�Ѹ[��fQ�=g��?q��q�=.>�Ul���Qa�'lS��;W4m���Jђ	��5b!KBK���P#��%m!O��B����u���ϱ!��0#�$���s7+d��Ѝ�`ِI�0o�G�����؜j��#Y҄sNH
��
�����LM���*�"��P*g�`�f~-<�Tu��Ѷ�T���X�1$A*�Ġ��1���?��������b�K��1c���
V�r����5\Dd�G�(��fC���~��d�^k��3�����R]'Y�z�y�U�Xc4P�����\�WN)#�<��8�N�O���_�dOxG���Ʊ�����1��?��Xr�UiH9�m�Z�u(n�p��ձA�U�m�s."않�� �����]��WeԲ`����I��؞�����E��oˆw{
�_�j��ӡ0����ET,<�H��p~
:՘J�4�K�̕x*�$�l�\�)߷��]�@�t<K�y|�i�sj<�d{�hp<��n��o�A��	�ӹ���ZŴ0��S��{H�g�����h�GV<�E�SB`��=�9��!���(���Bq�M��)��� �;䂟���e.z���
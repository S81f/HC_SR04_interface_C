��/  ��*pҥ�6��Y-�#p�\K���,���V6j�ј=%��K"��Q���>���T�mW8���GL���Q����LB53`��ݰ:ޫ�>�oa3�Z�&MU�i��êR���:�P;�F��C����/o=˴�����jV�7��eV���+��~+α^��P7&;��J;��2	9�3%��o��uB� !�f����ʺĠV<�0�D��<W�r\ǋХѥ����PPz]�I�:R��l�[l[Tl��ǲ�F*=��ar<��F���<5����#�A����2��V��K
�a�����P0m �J���rm_���"�;��H�2��t*f_�9i� �l������Ot� ő$�����p6+����R)�g��^���*����'���R⹛����r��G����}o�Y��P�&o�����3M��t���ai��3V��6�k����s����'X��8Ǿ��'�4{�
�o�j��g��U�)�J+_��M=:�a��|"AV�6Zvgԍ���]䢇iV��^�k�uDW��ø�Z#���'�I���E�_�k�p5L�q�"��R(8�ɵlcZBB������,U�F�F�l_?��a�#�=��IA?��{#��{eb�"��\y�c-�b�8+
����Hɦ�ER���+��؝|i��N�	>�[�|��@�f>s���AÍT�m�|qE�#�
>z�@s���K0bĺ#���(V���[Ů�H$��	��f�&d-D�'��~h_���Os���n�P�uI��"mp)v��:����#\Ox;J�鈗�~�P��c�؉�F�l�K���|n��LP�6F m�G!N��0%P�	pw��mD��CU��H2��O���%D� f� 5�U�I`5�.[Ëh8"c�����Ö�眷�@�o�ڰ����"�r'��$�V�p������;���C��õT(*�.l�?r����=4���o �b�I<8��ʺ��6��ڑ�3�m[<�۵iO30�u6���yI���}f��%��b4gh�ƻ�O�TyD��%x��i[e�,��\���{;�H�7�@�mm\@�KI���j�&PS�R����_�e�1���٦��Cއ�P��������a��7T�߉�k����룚�L̟�$��b��?����w6i3YO��c��Ӌ��r���M��H^0��ؘ�[�xYW���8tr]N��� B:�>#
�ʿ8�H _o���G4ğSm��u�5�P�y����U�G�VU\��U7�9fA��ʸ}������|���.��bXZ�p�ۈVH�g�A��4�RF�K:!HDH�����JDx��J��(���d��社����M<�=�e��tT������į��>>�4v1��p؄�MuC_��z~�g|�m��6�
F#��[������)w`64*�Uh����V�Y!��Q�A��4z0��MU�F �z�3�Z ����=�b��g��P�ѹt���2��� �
�m�O��]�K����(��|P-5,�?p~��a�T@��0潐u��b�@ c�Y�Q�<8�Fp\�f)iE��������x��,�s���Wm�:���
`=eh&���f�2�c_�� �5Z����Sd���JƦڔ��vJ��� <R4�1�sF��+V�=}�)���z:i�A�蝑�KA�`�������e�0�bGI�u&�RO��y'�{�5nD"�	��"�k������`p���9�N�H�r9��F2RAU#$u��b�_U{ܞ� �ʕm�6ĔX��/�B�3�o�����n�c��L�&=���!_�lya'��d�8BD��UG��V��e�ȧ�A�B=V��^�`�$z�%.���Eg�x�_M�G��+@Ue��T����E$O��F��n�F�~ƃ���FU����Y:�����3��"aJ�%DK��������G��K��z@��M%�c�v��a��Ł�?5����d�|[N)�6�옴�nO�uq$�+lu\`A��T����M�>�+�&!'����]�p�O���9�^4��XZA=�>�ԍs����BS�I�3�^�v	t+��s0���y+��y�2���cLŶ�4�w������p���.ͼX����}���WHRT.����~.ۍ=����e���Q(��,û͞sN�*��RtVE�N��@��\t�wQ�S��ǭl�]2H��	��NQ.]f�U���b㠲��_$�q��ڍ�y2tœ����ʪ�f"ur���)
�d 7h2���(��Gי�fB�3��
)�3O���62~�UJ$çխ���C�#�c:�r\~�V\�F��n�`
Ս�����]��.VAn~�A����'�����H���'i��ⰗI�n5����}B5m�Ui���#��tsD��_�?�����#�&�}jx�('LJ�:aH[�h	�V�1���>;��=��!�*�a�Mx� ���a�NG�dPl�B&�$จH@VXxk�eKV
I;/h�i-�3Xn���� ��6ʔI�� ��cD�7Qs���)"��6�1�/�/�z�a\��l���%��fzO.OI����4~������YMj��Ԥ���Z���; �#��^�V-[F���x^Q�T	S�ŵi.n�G2SFT��V�� ,���Z�?�d^���c��;��籾
��)'8���� +T�mb����ܯ�|��N��0GOF��_2O{g��i���� u�̩F�9��-��`Z�y���6��T�a�#^�~;ڶ�(	mģ����\s����,�:��/�<0�$'����O�ܝ�X�|��xJ�c�Șd�
Z�|n�n`2�5Ȣ/�R��bz�t��0,�بK���M�%�O�_��{>D���r̥B��Ƃ�~�_~��ZnJ���Ij��Z�cS��8q���Rz� j������,W6�0��V�%�fG'�^���ϑ�$���2@�7��«�x�"y�s=
���1@�3]����iFDh�IsJx�ٲ�}���=O�Z��Ց]~��!��Q�� �a.�J�q.͗�{t>�d+.k��S<��q���3ֹ5�ɣ-���P�����mV�a6s��=��J4k�Z��T�t1��w�(!��zu�9�ڒw�A9��aڳA��VEc�:mB,3y-�x����9���u	�5Ir4����E�a)������E�����"BAҏ���v��_���[`Ss��6��<�10\�=9H��H5�}6��=,=���<P�g�#:��񖜬Ô���Nr��tƔ��S��n�*�Ƅh~Wı=��MAF}IA���ňc��q�d�&-�J�'"�E�(Wf��Wӟ�o-��yM����t�We�vn����|���]��<	L���
w�2g�3	8�U���-��W|2(�	"�$pp#e�zd�Ͽ
��I<m@����Mx5=���8(�L�r��?��A�6U�D�A�@����9��h�����:K��_�n#��Q�}���"����� �PH)jh �X  ���P�a��ĉ�.�xS�%0�1��oVD'6�Dt���	���,B��4�v.�CA}��J (=�Bt��_����xu\�(%�ݗ��9� ���%0��բ����dayF�[iN���ACg�[8	Ot�K��Z��5P^!QD �h���GԳ�6�B�^�A���	�]�F�q��}���C�}�ćr��]�f�������pb$A�%�`(��~-�_�9��l�.@o�kXc����Xa�Z	{��.�j�ƬR���GZo2��	3o���P���1�|����������a
�� Qq�� ԰��s[���+�2i&����L�=71�+U������G~^r�ոֶ�U��H��tp���͝t�$�m(<��A�ͨ���rĊ���Abz2��~�
>c�n�	�����輅y����|��;��]>��~+�
7�y��%� -�Lj^¿�x�	���� ��q���8�l̡U�H�,'lD,m������	�a��0�6؇8�N{�H�|5��|�|
����D��7/xl}�؞��}
�Z�3_ǿ�R�;
�q��g���_��m���g�W��.B�7,-Ï�Qbn+� �0�R�����c���5o��Pk�_�����J��ֺ%M�"���唔��5�nb}��a:�D�1��)����I_�f�i�	;* (��0���zc�I����HW1��#jD�P���ծ�Ql:FbO3��V1b����sMI�N��ճz���N�J	vQ�V����}��v�v����X=#U6N��P��*ߠ�=qY��Q��S�G��G83��^%����ws���U4��ǀ���~����SzSt�4��e�{ݜ��Bq5�KG
7��p�卹�{@$ӷ�Є�|�l��]��/.�l��Ϥrޅ;�VK(KЪ(~��6�����3mbHT(�jy�0��R��|3j�ñ�zј��aD�x���=o�Vo����¹���>[|���fh"��1�N�儥u�㰵y��=t�M�9�\��;�*�rJ�h�M9D�h�R��QH3��t��(��5ۖ��a�uɲ�<�/�S������߃s���Y&O�.��{��3@ElAw��(��Z��,E�k�E��= JwfJl6��&��Tv�q��I��M��ɹ������M�S�"���ոI�s1z[��P�M�U952�;!��������9�DC.ۻ=�\4�azZl�R�XcxL����~V�1��p��u+�'_�?�.�D�3j,� ���� �3V��{֪�F���Cw��?ý<�m
юa2�ո�lkT��� �L��%���֊����^����/�A��Ь�K���%�v����@0x'��ι������v���+�Q��5�H���S-��E�\��˛9���n
��p�k|�h�f�a�d��oB�C�[��Q7�/O����ۢ	W9�����^��<�9�{�����0�˫>���<���[,R��9)hY��-峁��7�/�t8B��%�|P	ٹ~Fy��C'���Q�x�n�Q�h��E_�o�LM�,&�:}�����i|�*J�}ķPo-ɻ6���ڎ�pu3�#9��k)%PE�A�>������ʁd'a?%�\�Vl�L��g¯B���QQ-�:)��P�r�Q��x��J>`zQpO� �T+q�F�A��,�2���򅯐��-���t�M�� �^�l���D�W1+�p�/riIY�K���F�"����c�G�=�N��@���M��JpӮF��B<a`5�2�_x$h�%�'="����6�%��Դr�Ϣ�^�;�p܏��~��}͜?�LB7���]F�>a��`��8� �� ��C6[����_��y�T�8��y�v p2߷	:Ԋ	�
<w�3g)�S���Ђ��B�!be[J��IV�]�J�%�@
Q�C���@� *s;88~$��1��h^��lOw��!=;8�A}�>�@հ+�77)�8Ay����>�u�2q��Z���D�� �rc`T?V������0�ݐ�ih���v��6��ͽ�z�^�p1��&�� 9Y�&�h���n�1v(���}wt0`26u1`,m@I7ľY0�h�M�.6)���.���o������	zu��>��Ѳ� ȶb�.;��\k�[����E���_70t�����ە�f�;q�Ο:I���g�E�c]6���?SG�*�����0@��n����z���;�c�������1.f� -q�S���&ꉠAZ��H~����ﺕ�DZ���S��rur�XT4��i&��!d~�c�gْt�B˓�x�nm��t?3�K�ݿ8��
E+��MD��>�#��+����Y΁IhW�â�>���^�
�?���t��1����������Sx$9[گ��U�l�����cf�X0�i����L~�Gy �~G�n�UgD�h���f�Lï[�o�(LX�x���*�[<�O�
�8ۆ'�T��=u��%>r� �}���z���x�L���e�Z�W���q#�|����Â4W���:+9�<_���Y:�����T�,q�S�˴w����}YÆc���h�����(�jr�}�M��Z�O��R��崰�@�'�������	�#��gh��,�X,�h��\"���ٓ�=�);�?��L�m�+m�D(}���l���Z�H �kr���Z�R��`*�7���hh��{�d�?LH+�d��m���=,kFkx���y��9๦ǚ�`�np��1٥���4�����y�Pyd�n�xt�U	?8� �&y�h�
z�JǪA���m'/<��(n��t���kӼ�o�H��Y��Tا/����c8�|�Gb�ge��t
��/  ���t\����h(u�;����u|q�ak�Ӷs�J������M��=�Ii�	T|}���\�pq��d|J"�n��1j�30��ڢ �@����)w�U�R�s�I��<;�
��\�xZ0�L�=g�Xl!`����L���u��X+}�ݩ�h4�*�> ��c>%$;��]�q��3p����.���\06D橧��@hH�U��QJ6eN��f�2;Al�͓�Ƥ�p�-�}Д�)U��U!����\tØ��}sz�.����2�ȴ�l H��8~�u�V��S���QA.��-Rӊ"�d7�_U���5����tOV��
t$y�yу��Y��������3kg��<g)��#ھ.4��G���-�<�G�r��*��p��-�/i��"��a�]b�N
��}]��������\J?��7�"�B��}>���p���e����X�f@x6AgT.������;ʯ���#Z�[i$����HK��J�-ѡO{j����4��!hA�es����O8ǯ�q�T�ٸ��Q	�U�������a#p�طS���9�r�^�
�Z��K"�h&���F�O��$ц����s����S�f�����?�Sl� 9��G���X�Y4/Lǥ���p+u�fR1��i�lw��#�mȀ�n�p���2��^�X����8Ƴ
Q���.�k�׾���i�=*�__���V�*i�|y�ڀ/y;�6��8R�)�\��r��l�9�軈�I����'��ך�x~�B���+���~�e��"G�Isa+n�>0>b�4>�7����;�x#���������3&��x�|��h�+���	�y��X��0����6�ڙE��Z]�����>���"e�@�n��H�v��\��3������%��|��ƵbVE�F(k��i� �ST��t�|W{"l�8
N9�CG ��Y
�PI�o����Q���B�uç���9#K�(��!��,{>�R��>0�5�K�ߑ*a�HM%�J��i��<'CW�[�c�	��OZx�7u��/���#�Z�B���"?ha=���Af����C����-�����l��
��9�u��L0"���Q����ǭ���!1�n�}�"z�5.(�y*����~���z�p�<H�uC˸ML�vTm�1^�X����VR�~y��5��˘���ߴ<ߊG�{�ɑi�K)9������J�+��I	$����?H��џ8����}ɤk�`y�}�_�l_�FH�P2��]b��d�:^��Y>�_�B�zP�vW���)�$	7PE��Ү8�f�N,4�����]�oׄ�5�Y�I�s� �<�=M�I��� ��*jy�Em�N#�}���|L��Lr[�=7��	�ja���R�`^��Z�b����y2�π1��6�@"E	%�YJ�I�vzO4w<��\_E�S0����3(J�?,w���Edqz��7Q+��tfdhUP	�%<�JgJ���A*��H�SQS�$m�m��ɯ��(o���:�5�Λ
�����~���������r�6����YXI*�z�z� Uy ��4�x�x�0Ӭm�ƣ5��规ɭ�m`���Pp�͡u��
���Z,EO�g�8�"�/�0ܩ����sV�/�>y�V��J�����ʎM˅G[V���gN�[��n
hS��Y�%���۷<��(�cGwc���Q<�٭���A����X�|����@ڪ~�D*��,4ݛ��h��UWЁ��ɬ���cl���GذJ�l?�ɷy����Bg
E���B�3�FUTH͞�u��Q��#�����nd�-�9$`f$�4�X���݅9L����n�I]��sh�Bv��5����bw�@�LAxt4�����'��bXQ�iQ��Mf��y��Yr
y����v2#ma���Tx$3�ݟ�L�z%�m�n�v�/��dc/�EЀ�W�ո��Fi@������J���x;gޭP��Y�iLr��Ѽ�g��� 5}���8���ĨTH%sth>輝�x/j��{ɪ63x,�*-zމ�I!�\�$j>�%�F�axrrA9Y~�TcOR�c��������R�P��b��o�x�W`f|1�h�uE>�I����Ւ����i����&��U���sU؍@��$�xS��-��:�Wd�a$}��C�ԫ?��>�[�����C����F��&�e��{1R�b[p��9y�4�\���[#��L1�9 ���S.�w{/��%�84J��pw�L�)�[e�2��WT)����yS�7��|�T� i���7)W���Fs����s���:��G�z�b���j�S{'A�}$Eƽm��UL.Dyo+�c���ƶɲ }��,�[�ô :����m���x��6ƄBi��'�9�}7y�n���W9h�9��!�u����Ӵ���X�f�$��n1L�Δ�:�F>�#l��ԃ($�I�t�rC!���]o2�~�|��2Wh^�k�FwX����4 =�������m��*6rO{ؔ����?��9�C)g�9H����tuIJ�]*-�C玄 %��M$0����r�FK��W�y}�����ZK�V�q����g��	�	���Ƽx�f�D3*�<�/��p8_��,^�4��h.T��)HycWj��{��<dM#�kc�Uu��Ӹׂ�i��oH��2���ꝊĝLL��fW�^�qܷT<; PCLG���ާ�6-Ǭ,��f�(�/��EB���Փ����?�ʒ�&}�[G��0�z±�U^iZ c9p�Z�"���A����X�0��Zu�2����u��uQ�̋l>���4��hC�Z��9D�,P<�p����P50�ռ�h�Zp���WSV!���i��(n���U��Yʴ2
3!F�d�g"�<��KL����A�"T�&"�0�m!>xKT�,�6����]�7���5tP���ޘ��^��>�i^"���������'�D�_*jq�/=F�
��G#��%���2p����� ���_��Mp̸�G"ۚ�[O��JC0E
a�O,�j����s��T��r��b��B\G��ڝ6f�]��gS��\.���]�y?f3�4$K�^�x;��d��&ձy��r�YZؔp��]ď�	]���0��J��I�9�Ǉ
L�lO�_
!�yu#2���߶�"|CIU��x�]������	,VN{?,�+��3o��~<ݿYs�c��Ƃ��)�pc�g�Q��BmE��hõM}�-��:��z#��s���.��tNegyW^�D��,�c��<�P+F�~w�]�PH��H�� %��xa?�L;ȋ�B�h�������ԅ���{�@��/g�G��FbKG�C��ynx��h��L��R��^Q��N
m�>�A����(���?�"L�c���cH���#�4��5�=c��\�h�����@����)s.g+�`y^�&B��� Mʓk�w������K���[�^Ă��d���~Xl�%�\H�@>s_`���-B��q/�Lք������(=�{�S�o5V	�=�p����ɻ�@�P3S@}��K�y�T3�%�6Z�Yyw`)~}K���lV��BO�خF��u��;��Z��E�dX�%�FCBL6�Z��0�05S�Xg�au�US>�����Z��i@X�Ԋ���o57@�8��F�t����)���QT�-��[ٕğ5£��y�@��j��������.]0�i-��I~�W��:�4�_�	�����] �-*X����1��Đ�h�f���ڇk�ȕe�b������/6*��T���]w'&�[����W2�=X���`F��(6�ŀ>j�|_�{������ʨ�0Ո��@�a��5&�*����B��6gE�Xd�O<Y2������gr�_����8�j�N��H�ܘU�� @V1��ô�uYj?�WA�� �e,s��쎌�R����ڴv&���4�Z>�.��h;ނN,h��-���nY3��t>��ϣ&�iߥO;����'o�l;����"�v"���f��_U�th������R�����QE�#�E|�s���v��s�Rv�1�{�㩤&u��ū�6��P�M�؊���� ��`�lu�{r����JÀ��tnЪ��m�=^V����[�QՖ?����|�s����rR�SXdh�~�8��v��ם0�*R�	�!K�5�{�`�輻���0FLԴ���
��=��/r�E�+���p;��u).�/=J��ͷ(�R��:)	�JџTZ��*����z�=����a��1D ��!m�uA?��������|�J"��KJ��ꓯ2��'�I�=Qd���7�&���>q�ԕ	EO�jbԤ���v
/�>&:.?4Ni�J��`�*��r���_��v�N�;�Xi 	ZQP������_e�5�ƫ�n���+�WxJ��8KU��Q)9#
Z0Od_G��,��}t,z��|qhn?��q�d�\"�V�S�&YZq@�:��P�%�]�h���0���K�=�x�������X�͊#tރ,�v{2q�gOn�a��`�����A6���(�[��N�ݗ�*0b�Ä0K��c��A�>�ՒJ��E�V�W��pr�q�S�6��c�I����LǗ6�Ue�/������8X��I��SA�(��d3S�w�H�7���x����퓧(7}����A�M��$���`���,.OnE� �q��`mU2�������J㺐^�o�qG0+���m�؞ ���?5<gq �I,���b&�ʇ]9Q�o�˟�H'��80���k�<LW�fb�|��R�i'C5e+��k�q,�1VN�����')>��C���l���f k�[`K����w���.�FH�N ���<7�v���@ߘ��:.�S(��*�6 z� Œ����z�x��d��k��E:>�"�ƓY�kJ$�)�Y#��ʈ�n<'q)�=�[�h�
'm��` �eQzE��
��D	Z��§d�)E�ע�#�� ���-O6��5�b׃M�z�V��k��g�mȉ_�d�X�
T��;�3ƛOJ%tX�ެ��L<��W�I�=l� d��w\�5$��g���э���ό��c��@P�e�t�.v{p 4[X��oKr�{���e�{�49�7D� �@�>�����LW|��UNQK��8�.���H�R����Ѭ���i���8�{d���-�}�G���*�R/�Ifڰ@xq�N��L��Y��L�sɜTa��1}x���=_v�?�0���T�č�[�]|�x`�ex���,�ݷ|wJ�Y@oS���}ߌG�!��y�S�4��*��ǜ����u��dC.��S��X��v�س�˛���=�º��;�t�,ی��עOD���pjdQ����2O2 C<A���YEU�a����'�O��R�o3�Sr��� �U&4���C������5�^�����}��h��:񄧰�'�K��B�2r
tE��
YId��-�L�j�,k��O��x�/������+����T���vG���!h��$��k���.����Xܚ3g7IGg�)+���4�2CTY�Jl����~�� nALV�C�s�U�6>��{��;�v��VC����A�䎳�櫺k���L�C��������J�[z�Z{+H�hs�QFi���8�L���x�N��[�*L�%�.���MtC�5��LRۼ@�;��Š���/����3>j������v�k��y7A1��)�;�g������f􀍿��"��13�N�+'�=��Հc�D>��$��~I?4j���ƨO�.�����P@ǵ٘O���7@3�	��&n~��_��M��wȭ���Q������H	��g|q ��4�r�8?�l@�NIl��e�`��]�r��ɧ4�3Y4^�x���*�y,��+j�ҽ��T,�UQx�1�0	�
��������+&���S��ю!� 	5�,#�0����̏�@�x4)��H*��.�Tn��O��S�󚥸#�FW�F���.`�_�� cn���F��-�<Vr��ܪ���J���#K-�V���=<�9v�0��tظ��vOHp�h��!�W�+^��� ����%��"J�U`�x�bΘI&�Q\�Φ�r0¬-��� ������[�Hjx�z���P���`F��f&{7�e�t��&F	�}4���
fa����n�����1��M��${ff�gn�R
��0nd"�^E� ��1���R�OB��@���+�[�?�#�̘ۼ*I�SC���׳��S�>KVڠ��45
�i
���A��ة|�Z�Ҽ��Hؐ��1���#K
=���7�BɟY4ݎAD�)ܩ~[p�h��hӶ�������ۚ��TU� ���X�"�}�x���s" E�D�Go��|���@�AE�� F�0	�eu�-���1���K�5|)��(l�u�Q��!���X������G	�t����;�+�f~6>ǡ�b$b�p���o(��~���c�{h�_,첮�J�D���^�<��!�%��Ԛ7"�� 9�6��$@�U�oj�űL"l���q(�p}y6i�x��W���I$���%���o�dY9���

�z��w���i�A���$����´C���ΐW[&7�&�gĸc�͔2J��O��H�]!� >��4%O�<fz?=v̀@��ᓡqJ�}�+N2>�-.���wۺ�6%Qku#^[����I�N���d��n������!~'��{���7�CUQw���#�fa�T��pc�X�j�����׎4�hE'Cn��6	�?������g0a4I�*S�~9e�)?0���؍ǐu1<�d� ���-���y(�I����k���󽲫�L-��S}Y�E!1XJ۩Uf�`F2>*E1���-�e�#��E�g̍|�.�t
9�%����W�ր�h20O���^��Y|�A/��̌H�<��s|�վʎe�"�<��0A��u���#V9����Q.���k@w"ѳ�x��K�����x&3�Y��\��e��_�k�f���a��b&�200T�[.kx�Z�cA\�)��;��x�J��\�0��rP�}�g��[�_��U��}	�@��@�j�,>w��	oB�ۈ����X��s�R霺9�1ad�Vx#���0��?fF����mś��έo���슷]2Ʃ��e#�/+�1V0�ș���Fd�'0}���˫+��:2�"�`����|��a�����L���Q8�۽�7���,��ϸ�XN��R��r
O;�#=�X=oҒN��7�I(��\���'�&�Ī�9�ɯV+����S��̷�����0r� �+Y���ځr~V`��V�O2��h�h:|��e�ͬ�[�f�?v(k���/��$pZp�O�
���ƌ��R&tL�sl��C)n�}Ցs��fϗٳi7 � {��u\$��\��3c�����"飥Y���ځ&�"_����쐝�Y��b/��d��)O�}:�U�i���"~q�߃&���2�re�
0�@Uu)L����8E�Qp�//G�n(¼��ǶO$ۇb\����=��*e��^#��`�葦:T���l��K?�t��Os��aQ�v�@?k��0B��cA4Zuf����}�����lJ�l���UbC��1���~-8���Z��&@�v�r#	:���o�{�*���O�_��%��P����SD����L&"�A2}�z7k��I/.w�����No3V�&H�1��S`.q�H��C� ����q�n�Q���ʩ:t���UƯ��:�ګ�aZ�7����+����״�c�T�܎F�sP��3�Ҍ����ro?���ɇ�	,��4���@x>�b�W�O�z�WY����w��P"6���o�J"�����u{����pc���[�"<+io�G�t!�r��:�V#�-���row2��Lvo�����2��t_}�+��Qz�)qR���k�p2%dt0��Z�f!��򛳭�0��d�~��ΤA�yBz�M�`�J����� �/>摁�c�x@����F����E��
5����r�������O���ɜ3Y��Xd�0�Z����a�Z��!�}��@�h��V�Z�G2g�e�p�fYύ�&l����ix\��;��"�)+y3�>�mभ��j�F`d�0������DT�ـ爿7k�~��~e-��Oe��P��4n�����D�26�r�Z&i_��t� O`�t_�#�.-<�m�@��!`EY�{yS_��NuA*r�[�&���Hx����] w�TU�Ds=��\�+��4������2�n�껩����C�ۻ앴��Eu��=�+:e*�8�P] Vz��yO��2�Zh�1�t�7:ڭ�N'X�7��;�N�C��I4F���/�ܨ�~]�����\dAwX�N��n
�9�y�@`�>�2��Y�5���"W�R�iUa+��)��y�	��:e�Z���a<�5]��4�Z�8��������u	���pa�#���ō����/��V�W��;��q-�u�D¼&'26�JB�Oԕ�#��.�C닃:�3k�QC��um0�X�um֢�&�3��)��4Kq�A��K�&C�S���;P�r|��ً��D�*��\g¶h\j�E�H�2TU�H /�|W�����E�Y��b�k&x�B,��FCF��Z�;�CS�B���]��K��p}��z����,;ќ�^��"SdtZ$;�޸޾ls���X�G�����f�!�>©����w��>��)%���"�N��}y��]�N��AŞ���'��瑭
a�×��оJ���W_�3~wp+xS�#�*bB���c�h)?�+�,�G�ep�}��%�d�`���t�����WtO�ɶ�w����>�U�(��-vT���y�|�C����E�k*�fF\iR�+���M�k=g&3�;�.�� n�'O��{A�M'�;��O͵0=B!��J�Q�V0aQ"������2�2�?�lUp�<�2b�М���A�&¹�M��q:	�fb�'���`����%��'�C��Ca���J�3�ԭ�5��n}n���Et�	"�YSJ�z�v3ha��s�[J短D���𕸽�.���捬ʻ%����t�������Z;Ne��O^O��O\o!fcM�b��o	��8��Uڴ�ӣ��25��L���އjshb6��\��*W�k|�<�%�w������ /��L������;p�q@���q���8w]�x�jȎ�[���?TG�+��7	Qځ����ܘH�����;�e)]�"]k?���1?������m�k� ��L(("���/A��i_�h�Z,�te��Q,0���e~�(KX��lm���־2��
��ML�%K�%ڡA�1Ŕ�ˎ]C��������T���okF�;֎���hz��lv�T�Fp:楤���`�Q���n�hW�
�Y'�6]p�B�v�� S��}����)�[z�v�<�}���1���r:֧�t�!	�x�3�ʲh��Hzb�[�A6����-M ����Te��+�J������¬U�l�b"_��غ.��#Q"�s��$�P�k��j��P� ���\�7GT��d��@��ƪ�{#?z�U�ǭ�g"���K��/� �~�؋z2k��'[�dh\�X������*��6Z=$5�F%�J����;i�X��C5�H��zE��0 ��� ��l���DF�YI��[�j@8	��S/j戲C�`��rk�7C�!"��x	O/PF�{�$��bɴ讫R�eUV�,��;ڪ�x��]R�5�T�R�kWSR�����SG�y�8�)[yU��;��f30�O��ޟ�'ˑƎ�6E���b{>���_� �*0MB`'�@�K?I�����ew^j)��;���m~"���ET���T�ի`I�G���	C�?_���-GOV@�F!o�}A��p ښ����`�fR����
9ǱiЖ<o���@�^��B��e�[�W��iݳ�q��SB�L��'���i�,B(��n��%�L�9�Їٙ�0�c���󑹪2��>���%���-��-�G����>�#U�L���u�,]�
k�J�'wǡ�Ri�S3_�p��jc<��̀Ɏ�^�}�G�HK���Um��2*�t*�����R�፯b߬����������a�K�uQ
l]}.) O� ���n
�!%�=��(���{I�1
õ~S_�
T���G�W=�Z�l�[���y�����M�ż�	ZI��`H�5�$*��ޗQ�(��-������cR�E�f�c�I��u���syh?7Ž��)�҅��$���$c��)'��K�x;���Q��ͼ���RrB���*��Ce�"S��<�'|fVx��. ��R�g0� A*�?�y�raf�]Lq�zd{+��\���wF�uශ>�mW:I��h_���4$���P�=��W�<���;���-�Φ�6ձ�qي��誔�S���c���������M���O���l?�� ��~�n�4!t5��ξ�V��N�j�>���EI��`��ɔ�An�5C5����ŋ��`}��N�u{��ִ��3n�5i��W�1�2�O��A?����2���7����׳@m����L�b!���nz�iϯ7z��oe}RG.�s�S�cKg6���5h5�ۻ5�����\�2�L$G��2��SjM�FSU�,�|-�� d�pj�K5�Y�������/��?�S!��}�)-���mL�F�d�~G0�'�;�z��%=ʪ#%Tz�S�V�ŒiY,�N��-�1�f4B`��`��NP�i'�u�Q�8���{�-TMo�d��2���/LQJ�
H�!ٔg]��6�*ˤ����qѐ/.� g2}&�EH9��˫�{�b�Ab����xΠ0�;9nU��@��5vl����T&��gٚ�+t����!Z�����]uA��֥B�"���V��S3Zþ�Ǒ-1��
f]�P@=J�� ���z!":t��_��X|�~J��H�x�ey��\"u;��G:%N}����8pV��.3�<�mɆ�9�r�J��V7��I�l���w8w�%ێ���ք�m�,ײE���P�C�wjnR)����f���ϑ#��~;~�T�
�y����C3 ��u���͂5_pi$�]� Լnю�� x
S���Z-� �_+wx7�7���n����;u��1<�UL.}�I�����Z��G)�R��^�./e�"��� hV��}u�e��k`LI�dgKc%԰0G�݃�anr�嚼��糚	�J����g4��*lܶt�,V/V��n�撰f+p@#C�y�Ő��-�1g�ЁX�E�cp�-��Xd�(7�h�˟K��Lq���}oP�?�D�T	2�����]�q��x# 3���rРO�B����B�H�)�;���Y'�D��`���W�t>��'��.��"�t%�l�c���p36D�<cc�ZH]���?_r2�����D�.���XC���3':��f�I�����l�	9]��&��`��� �5d��ԇ[����\���8CK����d�U�x��+�K��ټ�J���^M x�E��ܳ��^v��l���ـAsU"iip	���
r���
4��P7'hzBX�R�f��;�}�a�[9�P�>��ٹ��w!Ӗ�)��Χ���r�x�{�=��,�Uѩ�4MY9iV�֠��²��r ;�G����&ͦ	F�^}�-�tl*घ
�B��-�j� W�h(862�kua�hs�$�)��������ڞk{ v}�b�ř�^J��܁�5Y="�/�B���ڄ�NҞ�F�7�ә�	.��L9r�.{ڀD�8�%�C���b�zg�Y�m��8Y�@[k��ե�Rq4)��	0����ѥ��|��xR��
q�*�-�j�'4�X��3��i\��JHZ�8k�Z��E1���O~q��D��B��Mr� ����������#LD�g�0���	mP����qzȦv��D@���vG�n��|N,�Qp�-�ٜB��������-�^�����]l��:\Ӝ�
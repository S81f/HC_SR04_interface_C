��/  G�������z������F��� m��7ў1�F)�'����p/@�����Q���F��p݆�:�B�m̏�sf���	=.7��$nٞ(3��l4�ߛJ��E��<_}<bW�N�!xoL0��E7r�DPȟ�b��A�ŀ��R8ꪭ��h4�*�> ��c>%$;��]�q��3p����.���\06D橧��@hH�U��QJ6eN��f�2;Al�͓�Ƥ�p�-�}Д�)U��U!����\tØ��}sz�.����2�ȴ�l H��8~�u�V��S���QA.��-Rӊ"�d7�_U���5-i{��v@(*6�AƾQ��5��qߧ����@1 |��s=��������R�VS-~���L��g>�Sy�_b�dLp%��o�FD/>�ԇ���pk2mGn.*d�l� ?ߗ
�؀�>Q���0݀�Ek0�B�>���$I��O�&	���2�89�;k-���s�iև�z��"��A�y&�=���mK���@KbCT�5�=���x�i��&NՎ�л�Si*b���n�	pq��|*lE<o��P�2;��,��Qs`��r�۹[�j���D��c/��CŖ��/�����[`%`q�+��}n�1�B� K$$q{�^fa�o���5�(�}s:� h-.�:��n�:u��@ڸ=���kVxP�xH���~��q��ǫz1]҃{e�ΣG-]K���H�6�޺KEc4h/[n�0A N�NȊջ��wΡ{�d���Bh1؇�隣�B;x3��ǚ�O��/@���E��>�w��~�6��Z2 197�qh�����Fc�>�$b�)�����F5�:k�h��#$�۪�'L}	�XʺSLo.����	;e�3���?��[�"�(@3RDZ#!�1l��3�(�>�0d���}��) ������f�d�9BW�|�3�ri*zNO�hF�?�'��%���q��!�Q=����QCq��E�nC�8m��s�IM`,��o!�%˱�Q�`xO zBU�!n]�a����]/�a�b˝�[a���a���q���(�@ti0G�Ņɰ�]'��T��&�.�X
cY�u�!����8��X�1P3���>����8���\�L�2nG�{m�{_u͟���ѝn�?ϭm,m��p��X�^��zv�c������{�7x�)�]��Z_���&�ľ^e�{.U�C��ؼ����2|P�e�T��LE�@~��^�v�u�L�l$gܻDgD2�,ZZ��ǣ�/hY#H�ՔcT)���p�l�1j���t������=(<�ְJ�̭���qR�yS��r��L�_z}-��>�S�EӶ��p9HdtL�mر�4#�w�/�t�^���Ck��i��пB��B�.E}���FR�L\S"�oI�叹���1����꒔/dCަx6�Fܩ���j�<�@���-�Ci�Z���&c.�(a��H���j����û�1Aa97��F�=CK&-�#8�22ZX��NMva��X��i���>ڷ��/��h��S"�ʌ1��?w�Cb��Dy��k�'��p2o�
�����jk_�h@�H� T����KO���V�C���ٚĉ��il���O�?��|��RX�f|Vݗ�X�[���j�4��7��ˉ;Rl���h<���;��̅��\��}�?ξ=��x����Gd,f�m�|�(2-��O3a��䳿n� ���r��y����;3Oé��4����d�o�n�Bo<3�j��u
Y�T���P0�$ @��XF���B)ɼy��BAʃ�Y<4���,c�m�f�:#�Cjm��Q��&
T��M�����WY9�����b���J	��'�S�
&ّAޓ��N���H�N���B5�:��é����+�{����(�.���n�Q#�;��?L�@�GS����C�iV�E� {?X~bF��O��쉪��B�zȭ� "��逤��R�6!�(�M��D	+}����M�\��o�8��M�.N��B`�{�B���?����zw����ƨO,��q�
ʚ�}}^���2Rx8?fOxq��e�_)�yF�w�p,�Z�a�qm}<{�� 6����A�ˮ�xysg����d��8~�S3���QY��2	9�ซ��!��F����XT⍱;�J�F��\(��ٸ�<u;�D]�`��~�����L�]H��X#�t��^u:݋��z������kPJ�����e�M6�j��"%_��!��ܑh�4K֊L�0�&G�G�?��C��W���-�ݍ8��a�	��b�LG���r�}��=��/�Dl����ܕY���a)-D�i�҄��@�YW����s�:G������t����"����3B�1�x��{6����I����j5bo��f�?>k��2�I]��Ķ[�`�d�wj� �],���:AQvRy^&K�m{ ~�u=09O7�'"`Ҽ}H��������}~�x�4�h�2���Rҹ��^�Cw�0b�V=��ذ}�{�3���dʇ��Ǐ�1k�︗�pK��}����-�<ʓ[�x<��t�sW=f(��= 3L<`;�'Pt��V�pû��e�Z����U�{q�������?�ORG��Js�&PM��M���8b|��G����-�O�գ��6�0g6�K{u���w><eU�_�e�Ǖ<s�%iᑺl���N`
X)M��8Y0�rN&�UF�����X[P�q�?�2�z�C�7�!U�oJH���sʫ'�&������P��ϻ`uƧ��Z�d� �å���-�d�w���Φ>���ߜ�~W�Ba�J<�&0�!�b\�.>͓����|��a'�l�\Xw��JFVyx�9��0�s���_���r��0	��ѯ�+Y\���i�I(t����R6p	�<|K|/��\wy"kߥ��_��ܘ��J~%5������-? N0^��#I+�բ��������!)�bb!�jW
ë ��f��wa��*�nk�2�w�m�p��E�
���H��`UH���i�Y��1������0�-/V�e8�v��ntWM_
Y�ɳ�i��*�Hq��[�Yc��5��1�;�"��eė[;Ǡ�y��6f��d������<�|P�����z	��
��+yeVth�%�_���S3 ��g�ҏ���̐�����I�p�1o,���r��!Nx�8t��"d�O��W�k8a>��
V�"Wu�`���h�C��~&A�Mdֺ���b�`���A��j�zԚ>[��^u%�6M����,*找����oB�K;S�EC���ث��グ.���}K�\�����h�n��Eȇ��c�~Z������@����z�pt�ʴ�j�� �M�F��V�a���VV;���Q��rpn_�D��s� C|���X���)������p�j)*D<O�����D���[?�r�m��W��mN4��hK���6P��85��v���B�f&7�a�\���3�dlK�/� bz�	Q��|v�6���F�6{tcS>��������0��i��a�pv$Y'�V�`��H�"0���H!j�P�\����VYfm�(P]xy(`�nߛ����*��['L�|�'>�z����z���"�4Mlu٠,V]�����#Xt�U1aI��k-P���(��r�(�0���\'��������YT����C\�`��O������A�fd蟟��Yߟ6�(�L��j0�l�4�z��]���սO ��$ԇY���a��:�t��%��h���c[�jX��mO������I����ü.ҟmj�h�2yX�	���:������G/�
�n�Π@��o*P{$�ևD����{^�8��wB���� ��$����O�Lm�b��S��	�����;s�hТ�����ڇzfZFCT��,x���0����F��|�>���,��y����1鴯	��*����ĕ����l|U���zPĴ|W�e� ����\_����<�)���%�Rx��:��a�r�����G��/�K���R�J�"XB3�p�&~5�����Z1��S �Z1SL�bhx<�8]Ftr�E����	A�0��� qNWn��4_��`=��d��Gj�$[���^����m�Q�x�5�f���;�Y������{�Գ��eH�IO�:5Ŗ�kQ�M�}��u���E�fl��e�<��M���{~<����!�ϕwha�1��+��D$4�h��莈���WR�T�=��5�F��ˬq)��`�Ғ?"�ٝ����	j�7�  �@|�n���*e���yD��?�y����e��!�?��sR2=�sE�c�͐0T�*K[A�:Q��&gQ�+��{W�������k��)���#^��s�T:���2�:��F�%&rh��w�y9��N���*���wK�[k���:�w��uiór[nJ:ܨ�<J����Y���t�έ�az�H��*��ƾJv����z�VN�nX9�2k�'������_�D�@c� �_b����4���DYh��N��G�R� ��E[������I]G'
�F�#�h]�8�:S2�GIv���]���8�+�R0���>_6�o��ݫ�z����FCcY1%�]���OT���Eɀ>��f�0;7�Z���1�/k���>���f_y����]�����1B�\��	q[ܴ`�I�&�._� n��� �����,� �C��־�	 d>�<��rc���pr��6T(�z�v^yH�2J���l�:\�9qWH�����w�����4�{5Η���t�+���8�av�¨���;�)G�n���jY�^�����_���dI��E�}%��{�(��N�%��~���A+�S�'"�U��_�Ҍf���\����~ŽRMC&��.]�gh�e?Dm�F���#frޙ �翀G�ca���\Z�������qjp�ӎ�hjP柏�N�"�Q��A�Y�w|��X�`v�>��n���W�|�r��t�=z9��t��ry�)��/m����R$u1����%���1l������cR����1�倿���Pǈ���wr�ؙ� ��� �el����⧲@�`�n���Y�ҿ���c�tk#m ��q�'W^�/J�4��n�>�M�	��H�4�w�J��1j�KG'0z�n���{��
�BZ:ZG��>�b8��%Ė������&����z�<7����Qlo�RF��EX�����3y����7�0<�y�d·v�s�;�U��L��GUZ�}����@j@7.-r\���?Q���k*4>T�G-�N�k��G6���xYvH+�¢o�:�qz��������ܪM��)�W�F�HM��0o�Յ���(�0���d���t�z��"kS� ߞQ�	\]�/E]3`(��u�=���m1�J�4�N.+�]a��c~_3�����ulM+/�>�uZK� ?�8�u>���oXD
4�8L�䱫���`��Em��-�V@�Z����v�����{\j�}�zK;��*4��Z[9��.������u]\$�1*�<�^Tޔ��s�]آK��j�ҿ�X�"D}�%ZGgu��E��x���O gGq����Y'��B'�Ja���C���Bfs�rt�Bp㙃KGrM�P��%��W�/[��M�[�'C�����\��̳��|e�G9@�7��Ϟ�5ple��:�zW:�
��<�����J�FȦQ��7Z�>&c֌�$��'K�죻C����.���2�d^/��r@�$>
;��Co?W�Ĝ���M6t��o���r��q�Z�`1�;�r�G��GP��{,��:��(PP�'QN,��f�����V�^�Kyj�=ha"Q4��j�^��A`�Ü�H��U/�eX��7[� ����8�Om������T���D�e��'� �/�i��p�_A���86L��İ`�ߙ����6h�:�8gH�����2��j�-�wk�c��d�$XBeӐ����ܖS>��	���BMfЖk��M$ɿ! d�I( ����^Y���6p��]1����xL9͖\7�@���	�|�^YQ(����0:8ɪ����L&uj͏xALP�_���-n7���% ^��ȟ-�!D����������ޕ��a�q=��r�0��Bʊ1Q��3�'籸Z��d����39V�q~l� BY��@�����(�f~>��%���KXw48��c��,�+W��1Z튩-��uՀa_��Q��<�=����9�0��E%̸:57�����"��ی���x��L�N6e.�Dd�3�HS�06<g���\)}��횗�lWiK4��Z��@j֙<��`���1|��|ܙ���Y[�'M�R�F�?/�:��C��U'��-i���@���)db�1LNXQ� �	^� '1�(B���L|2�X��ԭ�N��]2d���ѷ��7�3f��Ҩ@�zݠ�lM��H?r����o�?#o|�b['�mJY���}�;�Ïr�<��:%��Az�C��qe�P�jhsɻP��/\e��]޴�2d}¸�����_����0��O��}��;#�E5��ry��{�o�>��qc,��29���C���L.~m�ע�)��1P��'�Kc:�ə7p_��G�*k&�2���܎/ u��r��p��p||(i���~n_x��s=�5!}�k6,D[r6�>Z��m��x���Z��P��i��؅����AA=�4_���ωK�`O!�a��-��d#ѹ��;�'In�����-�N ��|�]����rΕ=r%��ЬEad�}lU�;3��vL��Ԫ��Nc����%k���
� �F�%�	���F�bGG���U������X�BS\��	��2������,x�XNרכ�ʹ�ܓ�R����,B��fs��d_�'��i��CJ��p�6��Rh�9��M�12��H���c}�6�}��ͭ�IT�ϐ�v��,��v����`���.��G���D�7\*�"��V���0c1��3�~�$Ma�8/�O�҉������d�-��(�H�p�u�8�ʛ��5���[���{Y*O��P`�]��xN�C!�|c�wB`k���)�;Y=`���d%SV�P�W*���+��aw�����Gѧ�I���%�xߚ��uO#[�5A�?!�������Lr{��鿣��	kQ�"g�k��4��az�J�(@Z�\��b�5�y�W�����!w~*��Oࠉ���Ǯ�J��ŵDҁI���>͒��P[��Q�ĢY�fc2�R>����L?�&�˺_���2���5]��:�=)+{-�ӉF/��,̹&V�)0�d/�`�Ƃ������5^��D�T
"��0�ɔ#�Ư�o�R�E1�n@,�h$�tth�U0�Łͧ	��>?㳍�Br��1��AwS�#{?�V�]l����f��J�JK���[h�!��?��9�����bah{����x��qI#��FN�!�Vg(_<�֍n�G��+��o����m� ��$�&>E�ރ��QWxLlG�t���>�s�'i��˧�@S���Jvx����J����9�/��P��<���t�af��ův��6Wɳ�|4>J~Ԩ|� �M�Ȥ
Zu"kNd���
��lR�r�[;ȺȶexN@��>��bL����6=�d��$�dsn("S�ꀋ:�/�M���D���G�;��U��^Dux����x7��:%j3�0��Co��j��}"�0Z�DK�[��ͪI\������8��˃��z(��38��X=
?�6�m��&1E�D���-�[2oJ�"0V����h��r?�@����(��!��M��yp����K���,���p��;��Q���?� �p �i
��g�r�r��4(��t+�0{�r���R
>�p͆U!�u�O��w'��mf1?;�`Cd�;�nl!��+�-ƽH�Hu��C-��<b���ȋ��y=�,`���9�}_�BG�>�(5N}]N��C0�	/~=���S�~��Y�u��e$l*ٿ��mh�%f6�; `fT��f]��p���t�1�����<�i��bXo͹0qA�b�%`�Wz����Ń�$@�K��x�ͮ�=GË�C����[}�x��s9l��ԫ_R�f����k���C\��6�� >p��R���	p���抩��4e�Z!�`mY�����$����#�-XBlV�[4s���!.PɈk��^�q���*[!L��=�-�=����DdB��{;ok4��v�ƒsL,j���W
ע�/��D��\K߃4oG�yo�Z��M'^�&�x_ݚ�YU�yq����*�^��`;=ֳ��u*����*��7׎��M9���%�
�=uN�YF�*./MF�̙��W�Fto�&�x�壣l d�}L	����-@˒�W�p[��@Y�u̧C}��Y�;�~LϿ`u�+����B�IaE!Y�>~�]`+�L߸T�Ee�X^�����*�LX����}���Ftz#.�Jޚ+��
x ���� Z��k�Xd�`�4p���Q���5TEE�f�E�k�p���*���ķo�����g����9P�%u���
e*�.Ǐ�ܮ�\�����3Tm�ꁾEa�cr����h��#��I�!@�S��C�Ф����q��;���/����3c1�pgS���R�#:�a6��|g�%w"�����Vn�t-�9ŕ?��^\��Ɍ��H�\WyI���V}�X:eدk+���c��� �i
�n���sg��c��@�4�y-�a�T�7	^�K�W�V �F
�6=>���Q.�OY�7������d���x��_����D8�S�a�)�Y��/	^k���L������.9ޕ�P��JѷĿ(�yju"V�����}),'S^�k�xC޴�k���~T�h+Z~�X��<M�x�R�_���	ctр�5��mV�o�߉P~ǎ�� 6����K�u��>C�P��;32g��~��k^�h'<�!�P��� z2�;irO:Ĝ��Ȓn�Q%5���z�!����)lJ:`��n!F��̅��ᑟ!�����9g.QE/��X�*e9X��	��j������'|��#d
��O0-&�u�1h.Q�0%�������QY���5�y����.V�ю����uѹ��W��2�^�ܴ�.^��329�<��v���ɹ���(i��9�۪�̶��]�e]b	�	��g�{K���0�l��5�W ר�Z�K�{ݫH�A��#��:Q�yGĮ(W�B�'��b�Jrt��8�7t�6ŧ���h<��s���F��T�>`bׄns�&r��2�U�e@�⎋4㜑�?�o��4#�P�o��� �m�؊r�l��v2����?��S_����iR\��*�k��+p��!|�"�6���'uD3�ކ�wbb*[v��m�nz�N'�3UA��d;Q��أ˧&�����n_���z��_,�R�����E�$aA�oXG�'zʖrpq	Ϸ�g6��r���S6�'�z"a�|+݅U�H��}h��?��LBa����1^q�u�1�=�m^N|Ս���a�����?��qs���$��ZX����ˇ�'9r���k��̈m�3E3>��g�Z /��3Qz���Ϭ;���nlCU��GO\t�ig��o��ϨӞ'�a�?�z2�>6޻0��!���.�Ks��h�*aF�+q��i�9�}�5O=P�� ��l��m�S���g�5H�1G�"�`��L�x0���K�{_��q޽�����|�*���H,r�n�C"�����4�b�;�mƑ�����^D~��'I���(�uD�\��I�{0P��oҔ���N,)��Z^s��T�灺A����X7AR9!ӱ^	�}��S!Ht����I�^m���&�ܻ\&M�-��Tr�0�4��#���Q��_��3��̋j�bsZl����	�枞�JR	 lC�s��0��x��*��v;fy���E�W�H�A�����Â.�
oR0�i٣��7�aa�Ϡ� v��l��H�.��SLo,�j`m�ф����fE)}�g-�K˽� x���\[Φ�f������B����>`O��PC��d�4|�П�8x/0$�I)؃�0�P=`�W�n�]�q�U�'=h|�4�X]ᚚ	b�+��e���a7�$oDU+������F�8���<�z�9���d�WĬ<��o9m�u5���@���7��I*��9�?=����W�@��֊�L�lVʿ������e�G/��k�9��g~g�� �rs�7eӵ]��H>��{�^:ؤ����K���bH�/Cd":Q��ǘ�#w��VB������R�ܣ�s�،<����܆�i*���<b��B��Eb�E��,�+);QU�	ʍ�N��L��_X��+��ʨ��o-L�iM��(����i�k��r>��֐��i�P��s�����|j�6���ʓ�S���ߓK=5�u�-�PK5Q�}%2�v�ZÁ�-u�,���=��Ҥǋ�)�Bb��-�]K 2w6.}d?&�K�wÕȧղ�#�F%�w�'𳪴��_S;.�n9{�ѿ��d#�e�Q�����n����85����LuG��/�ŀ�璚=.�a�@X-#���<�"������Pr��;2ӭ�-W��&�Ua�#r��9Y��rz����J>��86R��`M�:��D^��m[~,<��c
 ���#9�B撘������=����	��S1ɢ鈴6�֨�c��_�i$�ڀd$���/%���Ξ��Q�Y�5</T�Ŭ���_��n̉�>Nu�)t,�y�9��i���H���� �;X	t������R����7UA4���֤����F�sUKU/�������8��^�xڅ�������ު �Z�����~D��&��̀A;�����2�[���2>l����N����XD"� $��M�VK";�ōEl��>��G�H*U;&��������fG���A& F�����5九���'�F�{S
Q��~�g��SU(!��qӷ:P��3�eqQ�j&'9f�h�  �07<P���K�_�.I���J��\�<υp.g��S :x�,�$ d�`�X��*tq�`� ��W�ڀdq��2-@c���T����*/�^~/�(tB�<�,�ߟ�N�d_���Y���h])����\7���������+����e̗���O���U��i&:M%P\��hq	� 7�����￘P���z��X���~���X|�"u�_�d]�h{��,s����}�w�o��J���<��%���(O�[gM��ؖ�5�j��j"�'�qS�u�wȏ`�\�X�_zU�J�|��H<���;��9[*�B	.�3�+=goM�Q���|��1�R�^��x2������w%:A�y>;�Is`i��S�0�{ܑ��x�Wʦ[_�׈����l����$�7��_^:��L�s�^�m����/U��x34Qqt/��?i�'�K��7U��93U���$���ޟ�A~D(Y(�{쿳K�ӭ�p%�
�8�g�ju�%��(���$"a�V���$b�*��׿b\��G��˄�D�c�N�'�j'"$U<�6d�т|��%�9��j�(����U��Ol\�<�ז輗�vK�|F/E�3d���g��=�R�x��K����$?�/nKz3���pr�෣flq^�oQQ)��@�a�l'Pu�J�u�*E����V�i<��'l4�u���_t�T�!�3����]Ĺ�����&��qM3~��ڲ��`n�sr���;�{��I�)T��w Pr?�U퉮Q�
�%j
8�{E����@KV׀���ݒ�.�J��m�X/s������){)C��_$pu��(�O$�V�*����s���~w�h�GB�"͍GQ�\��.C3 �7���?����� 䳑d}�謊V��)�@�U�o8Dq�7�.u���F=���js�\	����J/�������N��ϲ������KvD���\�p>E2��n��E`��P@�	���za�1��W��A�$u�ڢqh @�a.g&0������n7w5�r��1�MbG
�5J�����mn�s�OdK��a?^q��ޞ~�%W�r�d�� PV�b�����L�i� V�$�rޮ�1�Ќ�HS*�狎�Y�%�0M�:��K.J�e��P�}�	�����URZVt1���}}�e�iKXЉ��m���`!��Jv�}N �x¦B;��<I�345��,m��ڀ����Y/��yu<�6P�>�sU���,���Q�h@��8����}�B��r��p�#A4��] �Ii	��x0����6:\�3��ǵ|57����Ŭh�K��)B�٧�2�pɞ�Y���e�l�������H
2�+J�zE�Ӂ��NQ�XU"p�5���:����1�씏+������\,�=�~��?!�~���3G�\��M���?^R	��		t|N+�����PJ�I�����IN���ߝ�7$p�+p��,��g'�e�gx�m�0~jk����,�Ձw�*L��G矁��M�(�4�h���<\rҏ���%��oJ�%K"���׵`]���Eݘ��>�?���+�����B��m�u�Y���Sm�N�J�"u����t�5��%R����~wF�'x_d�6t�Z�G6�>*7}t�����е���̩*T�UI�X�0�b��c�z�88{P��/��a��LDJ	�K�f6bh5���Hx�)B1,K��
o��4���H5ej�v�`�$���Y��+;T�
��6V~�I��8�~_���׾Ks�XE��,]�O*ϡ�~�y$��g�u�%�9@��#���0��Rď-���}]�z�f�,��<����s`�h*���l���{�h��4� �0Kҕ�Bր�(ƀ�����˨L �>}�k�R9�-{%a��>5���f�ۨ����X�\H����ᥦx9�6ʂgh�q����!wIGa�1ň8*�TXv�V�2{�ĺ�v(��{>��"ꁄ�^Y�����$[l/��?ݣ<$��ߛ�B%J}R#MOkʪy
�V�Rc��وkAu��Vo��Knu���*��~���t��=*l���C�������F�Y@hhj�bc��	N&�x����Q��R�+���B]�-u�2�w��$��,�@��}{����*����B�R!�(ye��Z.U��wf�`��l�4A^��n�Ovd�*䂯����c8w���n�k�b�f>k=aT�r�> =Z�A�~�-�U���85�U��g�H�fK�P���0Sz	�@m��_"��j����ޱ4%P������Sc9��R-���%/�q[$�R>9���%N�q8�1eRM�^���j�(4���3QA2�7��|�v�4Mr뼧��3�N�P�L&���˱T��j+"w��`��w����a5͒ޜ�y�˼n�"P?Lrɋ���+�kh��vHK�
�%�����΁�z+X���n�#�Y�C�q�K
*��i�ߧ~?_��*���v���%�������ٶ��L �Uc�iS��,N_���T k�:݇x,X*���4��E�SȢqˠ�(M}gX�@>ڑ�� �[�@���Bז�1�v'��@=l��`���䰼Vm�:�hp4���I�ޝ�L"%Ri����h�l?�W��Q)W�DcwtWh��)o�=�����/z
;I��$�f��:�<�$a����k��}+�"\tD���˗]��*�$+Y�7���a��u��G6'F��#l߃3��}��)OFz����S�VlΚ״�D ���9A �<c�8BP�EK�nY���r�$~�P�p�T�D���b6�IK
�0��YHa�rucbVK1�S��K�\\4eq�C	��)L������l��W��~8��n��厀.���smk��,�rhݢ8:F�h���_�y�ڤ��U9�~��݈���sQ�UrFU�K8�w]x:���O���lBHfY� $��3y]��׎x�T�
D�"&�|&լ�?�uV{�jYa.�x��N'	G#�G߭2�F`�cE�@z!u"g�W�~����)� ���qF��vp���:��_�^m�k��s��2�S�q�ɬ�y�m��U	�b���&C�^�Lz~�=y��nP���E�bg�G���|���"�
eF%L8�v���?A3�����Fi�������r�2g��H4��Kr*s�����3Ca��:��y�����u�EJ\_�m���4�⿕y�_���]M4%��շ�#xl��*����B����K�jb���Q�(���"\�H�^�ܯZFoA������V�(Һɋq�Kѐr
M���~4�H��"���|�$�7BUx7D[�wTG�/s����X�z��H|w�2������u�al*0>	�S��Ek��bX���2�n�v2Ё���0z�/`�i�M@l$,[>�7�C黭۬g �a�M�Q����H�41�8�� ���YXҋL��M#[/����������ȸb�[.�$q���U)���gGq��a���X��8Z�8|ɯ���T�����8��:��{�?��Fsִ�.$�ˠ�6%@6>o��k������K	"v��	v�V�=HG�Wo�!?ϴt!���ӽ��R?[1Ls�#�4��b�c�W$�	,.0��'�Ru5�+J>Wnl����8\�D�dzNP-;Ǜ
ƃFU}w�K�������!������q�8�,��/s�Ar��X���CM@>o5���eN:�Vj������6�o�0Ґ���L1�3\�]�8m��S^�������Z�&j�kfƐV��Kzl��o����Y�$��Q�@V����x��ep�n����ֈ���J�'���"��かu(���*�AX(UL�l�BfP9q��l��s旧����O�*��q�&�;N�r�M�?�;O�(X0߼��=ajG�Un
o�ud?�8V5������Z���3E�;�y�4B���2@֚��[/����T�2���30>рW"9(���Ɇ�L�@��f8����}�<��D��t�,�:�F���-���Wu�d%��y�&Wi����;,�S� �B:lM��#Dw댖�ݛB؇�n8���	�� �Nٵ̞��҂1�_Ӣ`_
j7�5A� ~�*6���R�w�Hj7��|&�IE��u��p�k�t~�@�!��rF��]�����$�߄NE����D���$?������g�	�e#m�VGhZ�{H����hFp��
��0a�6,�r��)���	�*9�޲�m!g7@���u]�G���@F�B���W9OA���b+���M\��ڛ�%20�gC^a�P(Q���ȅ��c7(�i�Uk��@�C�xA�A!F����	:������\��s0�ޮH���?	}=�~3�1I�B7�B���:c7n�L"V��t�ʛ�t{��X_����A֟'�#h� ��r�>��J���i�ϼ�������wӳrs�)o}⓾ą�d��<�&�:�75�nS���:�dKE�F)���.��?B%/V03a�cޓ���ɪ�O��}E�_�,[�f�ɖ�ڸ�{�m$	xP0\.I�j)�Hxb�-_E��X"4�I�EzR-*�{%�	��A���Ddo�W�A{�8؏a
��Vn^����������JAUr~L��-� �Vw�Iõ�5���K����N���l�;�-����qa>%�F����I�K�V�:�D�S��]SAoS��S����|�	��:��B�9�����jbxCJr���hXņ0�=70.5D#*1�/d3fK (N��E���5ц����bwx�S�ؿ�!oed���]+�wj@���;m!�Vv�zY�E�2��k��<��s���<�5�Չ}őQ�Qؑ�|�)	Bu9v�ݯ��N��y�2.�t�T�J��#���z��#���w��aj�A.j�@�d�S��~�)�qu��XOa��4�6��קQC1���g��<�$�1vƍ���;���L0qu�����^�fj8Uz���<�.?���zp:���m8�8��M2�g�-�~�0�ؼ�~���q���b΀n�2HMK�=]��l��A|�l�>������) �v�A��`��7oә|@�}^�\I��(�k��q�7�=5/<��&�Iy :���$Մ���7� j��*X�[ڣ�( qE���y\��t�t(������t	�ϙR�0:Tb�P�l�C���袣��{�[\��?�[%/"�k�`����@�c��*����Y�"�HVuQe�cv��γ؇@���iq�|�f�c�슣��=A6S^4㤡�dm����E��
1x��.Ę>G�9��Bw��0SyI�B@^=M`�~Kg�F̘�^U�!�O�t�s�^�z\�]���{��).y}�A(O�XR�������XWDu�ǣbOX� pO��ǣ��X�_+c�O�fJΑ��QE3��u%#� k�u�|7x���%غ�#<�an� ��i�\jH�N�/�y��A3�Xf�� ��*������z`&��Y��G�����B,����{�8g��&��t="���̛���8�wݥ�Y�J�^*���6��-/��[+<�+�XQ>�}�/V諕��!���F��H/�`���o_5���7���f���{'�^����U`�F�quz7�Ɗ3�	�эpT�s�S"^�H�&��B@��A�O��eי��<L�(�\� Z�&2���%�d11�p�T��22{�FB�3 T}|��24�Ű�HH���`�Eܴ�SUX#��.�_-�z��(]bLE�;A�ǘ��R���?�Ɍ�dK��s��R� ���'��9 ☮&2)N�')3�XOE�j��?���s=��(�#;l����{j��L>A2�m�]�QL�2BOtd��"����\DCu/�!fB��J���t��;@F��2�Ao��&��RUʀjt��71��]�Ŕa�H]q+��X��H�h|R��� ����x� ����uE!�|)�/��].��D&��#O�90'�׃�`;o�	�^��9�i�����K>DZM`���Y�l�d���Ű_�M���S���Rm0jd��T̴�й��Ö�͔�H^$��l���w� @�Iؼ��R�x~?���5kh��ZT��!L}�4�ι���K�i�	:��Q�O��<n{�j�:�"ִ�^���0�%��}ݍ_�r�BI<��TT(�����%����6P�قE�1�r�JaV}�N��^Xăaw/F
��/  #y��W��K�\��H5���H�=�������N�47Z�Tn���렙oq ����hgg%D�MБ��y;=.��i-�CIEO!W�:��m��M�&�{����e;#��a����LY�Z׷��qƲu.���� ?lf��.?�W�<�"�t�A*���u���h4�*�> ��c>%$;��]�q��3p����.���\06D橧��@hH�U��QJ6eN��f�2;Al�͓�Ƥ�p�-�}Д�)U��U!����\tØ��}sz�.����2�ȴ�l H��8~�u�V��S���QA.��-Rӊ"�d7�_U���5
������ݥ��?7�q���g�؎�J��`c�g�
*�:)aL�n>	aC�	[u�l���|^^ڿ�d"���M;<�&Y V���So��n��4��ЌQ\?�|IuƒLӫ�P���*W҇4�]F<����E-� ;���%і�2�4
���<�94
C��������B��)��N�w���#�T�����HKwE�ت����R���Qw0\5�7Qd�vͻf�{���������*a��h�%ϵf�I%�O�י�U�n%��Ǚ)e���V>X�G\	0V��1Z��"J��x�Z?�Y^nO�F�S�������axr9X��b��t���w����]�;b�ɹECX��鵘����8���"���z�T��O�&N0��?�G���+UH�`�]v�S��4:l��|�e��Ś���r��
���d��B�^�w����Q��i.'z�*��_R�Ce�v�'
�C�Tdꢮ'ot,Q�b�]_t3�4��A��[?��$&^
N���Ɣmy/�^3ѭS�1�&]\��;L�FfV�G�.C݊k~Ҍ<�T���ǎ��Jg1	�~]��sb)�%vc:F�h1>�La2nS��@�;��藲�`����/�9Qf#�[����4���\�,��̀�R�^�ϳ�cY>J����YWk�	��ЍHr�QyC��A闸.k�#)�f��xD�f�,�GY�rRƞB��p�Es	�f�]P~�_�F���[j����%��F�Y�����؉�+��@�G�o��f�"��A.�)Sʐ�ϳ�K��}���>X�:N����S�=��g�oN1v���P�8��Y��� �a7�^N���8(I���S(m|���L`�Q�E}w���Ns��"�mQ�0A'{���=�	p�vbo�_�H97zl���bj������tK	�B4�9��m��{�v�_恎l7G%�`Rm$l���jW���B�}4>�)2���s:1Z�-KP1��	-]?�j��@�73���B`�1�l�j�ѕ���5�^(���b�k^�I"#��<j��rfz��o��d�a|\�5���������1g�~�̠`}��?������LrI3Cۆ0��FJP�e������P|`v���X都Hi��`N6���F�]�h6�^��W���ү���ώ"T��$�C�"?��[8�E�����L:�q�cu�+d�"NHb8���v#�-��!.OF�j��R�]�JQf��ԕ[3c\����/���q�u�H{O ����ȸ����;������ǀ�m�e�7uʎ�e�~��u�1r�`l�s��?	r����6��E	�����#�2�0�A����d���VT��/XC�wg�}x� +Q�����F���&�2LN�A衬 ��G��찌IR�*�_�q󹸃%M�\=/게�М��f=hɪ�zEZ�'�_��v2(8�דO��ξ&�S}YJ�.x�y�|9L��Û�0x�+SK��ln�����|��P�WjF*y<��F,���1@�ΫSp���l!m�f�a\��[�%��t?���Y&?�{R�c	`D�1�.��E�Vlֶ��7��)��|&^���3�s`��p��%	��a�P�H��E���w޿�\������D���e��B�̀�0֏z� �1&���l��{���l&���lk��3l�<y��Y���"�K
B|L�jޤY�]��6����>��@�f|a�d���Ɓ��;�|�b����Ғ)�傫�ew1����F��⛰+`�z �I��� ̐t +��b��\���}}�|7�<c�s����UP��SAj��pl��p׆�r
�T��D�h]���t�B�d���=O��V]��o�mD��4 
�>��ú��d�!E�ޛ��qH߱0��I�0�����wT�q_�0��+Eg�����I+8r�����u�x
�$�^��3f���kć2=*��9A*�}T��_����B�z�5Q�+�N��O�y�`;1�C�g����
,�K�F5�V���︥~4�e-<�7d8y��`8	8�\f�2���<���q@���t��^���=v?K:�3'�ل��t֚0m�=��蟭�eWw����GEL.��\f���������������j�ΣѱCm�*�����S6�����Tk��dۓ�����/�m��Ba:Nc�,�ۀ9�0N���4\I}U��������9<���q	�=C��(Re�0	�;?�������t�rA���Ґ��>na8�so�Wx�1�*/(���:�B��g�W�`/T�����Y��7��ejζN����P�'��|q��>?�Nd~��T�^��߅�ٌ��͚�� j�z��Fi���\�mCݬ(�K���8i��L{�$�U�@���8�����`��ч�h��ľ��ޣtT��~��-�-u�H��pi����J��g�<o�M�r��ʗ$lN��	�VM������0X��)� �&ځ`.l���u3�}��,��4,���{x��cд\ݫ�.��*�8�R^����l���U�Zٴ�����E�#������'��WS�dG��n��G
��j�P�2�\������n1�bMw�H�ʾ�r~!���:b�Zj��58�G�vѻ�cQ"2)uQ*އZ��1�v��eI݋�Z�p���o�ާ�K�K�h�E�i���-��V�S�u)0��gX�"<J`�Z��S���@��!��NgEO�ԅw�����H�u>��nQQ0�9�W	g_��0O���IHb#�p���o�a���d�m���T�j
I!.�
lE���{�,:�HU��sw�*g��E�s�6�(��g�b�>�D�٫�H����
>����9�ߺ��/��7��H?&�]Ɖ:q��4��%E����=K2�2���5��w�n���!A�V^�U�M8=åŦ�V���o�|j0�=��z�K�<�t�u�q�s�5��54��a���mMy�=���)��м�
MI�3��be�V�%�ղ�C.��� E�tj%�-�3��_�H����7��9u|,j%�C�F.�m��_�G	we*Z=('�r�z^[J�I;@ٜn
+󟂄�p`�0�n��o���m�T��͌�M%7��Ë	0���I0*ܴ��ejQ���>7�������p�QX2-Y۱���G�����Ӓ���(͑%t@�T�✧2�u��a�1���孼�������{�:�1�ۢo{�'��	��k[&��+���{*q��S8mOҏ�;�}�v@XC5w�nBj��W�ոv�?�d����.�F,�ݸ�#����?�a.���	�+7`�c)�{{vE�Nl��eӀ�L�f)s�x�d/�s�=4�M�z�y&�]�Iy�����q4��K��q�O3g�+	F�(%�_�@�tǻ��sw�ً�߫j�ҟ��=B +��swE�����3j�!�)���ܞY��Ռ�y����(� 6?�Nv���l����N� *��Ɔ�dt�h:�A|�O�d�(ae��gRY��7�����c�V%4y�`�J�F(�e��"����W��R��}p;�)��	�e�N����w�h��ʄ>:�R��*�����%����Vy@̓���M�*
[Ҕ����,��� ���� g��0�Y)�d��sy�{�࡫��"kwi�v��Z�ݷґ�z��gzQK��BDi�MnR�H���htU�:oRdaժcd�(�c0� �VVl������HU�ہ�hwbEV3X�^�2
��K�1V]��u"�����V��cZޑu���>B]\T���锒lc�JIG�	4y��E:�5{OY	��a��Tgb#�C%���P6���C����g3�2OAӚ�K)X{L��u��?��"���1իF��F���H�6&ۅ7��s���T0�%���������b�t��Fos����7�,S>���+��ml�
�ѻ� ��,'r�=��Vo��-����:/j=a�^m���H͹�eEd'^5�� `�%����H���h��	&lث�~�����x�p~����3wv�ڞ��`#bJ.3A�5��q�HZp�`,��W�Ē��M�ǽ^�����/q}Z3�y�W8}�(���o�̍׫Z|;Pc����ӑ���o��`ǜ��d^�Cff�]pĦ��j����@ئYn;�(�:��m]H�9[�Ī�_5�+�/�@`�I�N�NO��.s�a���7^]��s 7�q��i��dWY���`�$�{ 4u@�(6��7[%B$�,�:���e�kAk�T?
�É@�Eg��y�ω���u�o�h�Д��P���'�����y5��翅=��Sp��t
�J�qH/6���C�<���Y����)R�}%�u�������]�F��&�D�~ER��Ċ�e��sv�w]�����o��o�M�Mb(��n���+/bӈ��
�S4�w���~��aE(Gî�/�vo-���J����Kφ��0���'~3��F��G�����h��h�kI.G�a���Ղ���xg�o�;f�6>���R�'f�/к\Yp��a3U���2L˟�?���g�Q*��9���V��HL��W� o�H�����c��:�.�#]�H;�4���Z�YH_�#�5�	�F7���p!j�hl��x�;�n3�����_z��o|���b��*&<���s|ov��'�*��J"h������:��B�j]D*s#G���y��9��`T�9��\y��e���+��4���c7׼���:~֋�L���Xv~5�ܶ��Z�X�mN���(�-�8P�C?��2����� ����T�y-H.]Љ�&��j��V����(������>�T��WS��93i�BI[נҠ�e�t�t܅00��D�{���*�_�� �_�Fj!*�Y�vj}�v)�e�����:�?D�����G�\7�?��˧iN�V�����a<\�쳹Z�O��4����
�G?&�p�-���%yg�	
��2��x�DB�8�۝k�6h	��u)��� �X�Q� @�"Y��:�C.`����}�> g����-Po. mD4� k���W)zR�*C��jńTxNn������_�*	����X�G0Ly��oSZ�Q�j=��3	�I>b�9��v��؉����>+��G9���!�u�6��b���?�����6b�� ������qQy�ȝ�$���m�1ܔ�^y������o?��z��Gt�t�8���퓤�a�unS���Y�F�Wuq�w�  ��IwB4�i�ޑ{�@8��MH�r���Mp����Oک[1�e�H���o�m��8�# [�ui;�*/P�Gh��a�u\Op�<\��p� *0��e_�OE'I���L/��X����z$麓-�
��&S�i�������ݺ�"*(����,�����6��M����R�'\f'��l&Q,b���A	���CQ���k�͘�"�є�����^ W�Y�=������Z�Tk.~r�W=#c4ov]S��ߴ� � O�FqI�n�c���f��������$��?j:�"�-�&Ŗ�iN��)̓e�WkD(��D@^�;wC�Z�ն���AG7�E#���֮��V��t�vZ���~�����c�|��U�����D��:��g n����mIU�_q�l���o\��Wq�T���������3\���W��t*\�2���6�!p`L'��Zs�#|�⫺Y,on�:��s"�n"����+4�iB ��"�S������.3Gs���.�L�Шq`�������*Ͳ�S	�����!�)0.,U^R��ݽ@v���ީq�lWų��*NɎmî�
�+�fSdI��Y`<�=����a���8m(n1�������g�Ģ�z^Cx�M����	����T������y�b��Y&]�
f�l�D���� ��Nѓ9�2�ϝm>yi,I�3���q�O҆��Sο8����N.���]	���LS��?sϭ;�jM]&�%�
���>�duoɴ��fF����b8A3j�V�2�� [��P�A M~��²vsm��	����[��}�q ��merQ-�F�A/�p���p��aԘBչF&�s��}R��rZ�����:�JJ),�������1e���ܟ,G=�<��z�È��D�|?s�ʎiy�� U!d�*�i��/܋��V#���$&��;#G���V:u'ݩ�!Gɮ44=���0 �
�"p�Y��zJ����K���[����?wZ�(�8�\']^I`�mp����M��^dO�B������L����*���Q�1��>�/�����u�
�9��̠_q�_����j�+%n�����z�u���a�B�����A����c�7]���M���eE���Y���~k�u�T~�����j(��)�*��u�/hl��W;��k�4
�?������}�r�
H�~�eLը�쮊*A���R�o���K޲%�}~ɬ�!������}kl�����5)����?����m�Ҏ�g��+����waU�!u����� ���Ů�~�����K}�+�}�ʙ��Љ��{����3����[ؗ(�9���	WThC�m�ٮ����P˥%�0d��O�,U���������ڐ��`���$^"���2��Sd\.�����?3�'6����'�@�K��\��Z5���Mߴ��@$'�%6�W��m��5��6�J&~L7���_��u��s�N�H�LIs��������r�i�b7���7f�4g�{�`�=���'O@O2|�z�q�q�ɪ�ǲ����<��m>8"�\(1��Ԙ[�&������Mp� a�Ԟa��l�� �<�����n�I���Xb7����e=Ks��9,��qǟ7W�M�	���#	w@ྻ��9E��h?d��+9��,+���>E�{�!� �V=n��RsE�|�c���}`���7"V��ݴ��!�m�r�4���/���-�P�=�r����d8b^�����A�W��)$1��@8NW��8N�t���`p��0�AU�dx����h�A2Q�:q���1�9��I@M-}C��X�͇ {�����)9���t�l�����軺_+�!eOT~0�B����V�K�� ��A�eŔ�;=�k�n�LA���XC��tX�Z�#;5�la����Ć!��y���7�}����&1�[b���"�$9�J;U|@FM��[����D�XI�k�((jW4�`&�Dp�<�/�~yi�N�XG�zy��y��R�ż��
��1�ո<�i�r�v��V�9�Z����v+�1��W��ɓ�kf��J��^���9er�@]yT{�S�N��s�٬6��Ko�Z<�7��k5��@	D�n^eL���!�A7{�د�"N ����Vy�2�V����75�+�(�h�gu�-�ɔ�&��!�O
g@�7A��ƒS�x�����=_ b�l%;�(�S�n7���t� �2��ˮ��F�d�������.o� �6�$Ө&GfH�C��_.Ntrn�Y�򹌱�k� �~���K{��A�h�"��ܡX�=U�����u���dK.���»����L���A������/5���L�� ~���3�ܫ��.�������n/�s�sd�=ŧ$��� �FN�=��=Gs�D���r��hF� �-֬��� �]�+��M�dm7Q�MG�Ma\�w̟yf)�wm�N�Ym�ܸ
�U�!�����{��Ll�=t�����»m9���"�'�=$�5�5qz���1��0ǻ�tL1s:�]\۷����a�A���hF�m9�ԭ�w�ׯ_�{8/�q�^��OI�Z�N+i�*f��,Ҧ����R>U�Q���!px�d�+��|3 ��rV�,R��j���uk����
�� Q��(��c��V�xӖ>`�m
Oj�JRvj�y�wy*32���<	�4�S��h9�B�~/�eyC����8Lt��X�/h+/%$�Ft7F��p���?@�O��z�t�k��|���)���lM� ������YlBj%Ip�Pуg�<�	��&���VW��	D`!�1Yp+���؏��N,�H�\{���|AD1祬����|d��W]��+�B�0Wy��
?PfC)�"�>�ѓX�;�?��$Z�`m%�(�Z���TF�Ν͚���������(s��ɲ�>�)89S���O����JY	�����d���iỳJ��JX���:��H�"G�������E�M뗦�R�o�Y�y�e��G+���ҩ	�1գ��Hl��y>
"T�bޓ8y»,
��f�K�xf�틳>����}�I]
~�q���'}S5��0	�?kOΗnlr�:ݘx+���W��y��[X_���|�����م{�*�1)�į��ǩq1��k?�󷓞�GH�Vn��(��[R�-	��O!�f����O��[F$�����M�T�pxi�l��A�9�/����Vp�wV`,lg`dgU�C�Er�y�����#0{͔8�K�:s��X�3����)/��e�86�7�"ڒ<�7
�"�M]�Vh��:HQ'����W�U�68�@�6.�]��JUעtIJY��]������ �^�5[�3������3�\�+,������^���/��\M#Ĝ,"���g�O���Z��R���������RU���<n��1��"�څ��e�v����9U�y�QTx���F�*��sB$�p�5Εj���CX�{zQ���C���E�h�.kvj�i꼎6������l���,Dǀ8����fiw�=ƨ���3P����A�ۏ5���Jn	�U���T�X~^/�k3ٽ��6U���s��W�Ц+��y\w��e�gtЗN�xul�8��iG�������F���%�2J�Q
���5z�G<�g�Dе�8޼DE�����$JE��W������Oe^�.C�;0$��1�琰�4fz+> Ť�5�1!���w0�#�/���@��Hu��	��t��a<�מ[��:���<����][����BQ?�[x|"�o�],��ݠא�g�.��rח\]ma/�9Ly1[)���*庽�M3B�.��6�V�[(��C��"�k,��������B)����om3���CLr�M9.'YG�&{ ���@�����}���3nÉ������w��/�8��Z��D��[��W�/A��7G��K���LRws�2��x��
��Y�3zޥ�\`u��F�aR����!g�~��+��!(����0@������I�lM�ru�m��I�2����r�	xCO�|�+��аZ�qɹ����8�,��l��R�u�A ���A�;H�n4
Հ�����3�%�@�*
mLh�E�}a�����Fe5:=�8����	�A��7B�M�M�K����; =N*
���v�����w7��1�笞������L\Sv�>����e)��4X�U��,�����; 3�G�q��{$���d "��t7ն^,x%��U�:��q��A�u �+Fbd*F���u�%y�S�<����7��U��w�{2�����n�alÀ�V��Ut�+����h��h��f6��Y��kT�]��⦭ �q�[$=iM��۳���5��Q�V���D�8��$���r�i�Ǒ�r�V9<HD��j��t-`E��F<\
%�4�t1Ǽy�k��@I��7md�Ug��P�9X*5��;Ggu��^	ºƓ�́�B��#1�)��ڭv[�F�*�G�*��xze���Dpyl��8r��?r�P�_V�2ؗ��h�vH��4:��Q����F�N+��X��(��j��<k�˞;�{�s�ޅ�v�|I;{���q;�724� P�	�"V�� Xy��Bd�����\�C�es>6;~��bW����x�3a�/�6z���Oܸŵ������v��.�tˎ��$ ^�::�bq��0񯆬�K<
���IW��)�S�	Ǝ�
�J�n�4wl�����K�ϙ�r�)R�4���\K��bS�p4I�,�:���Fm�j<tᢠ���!�.�����5�� |�^h��K��Hb�)T���
����Ԑ�D�����L��Y(�$VR:��]�^'�+g�����MiGXj�Z!jy~q#D���F6�A��-ٕv I\V����@�h"CFI��`�,�T��j�V���3(�2�0��{0I������y�X�	��<k@�"Ɛ��C��~F7j��b��t9�+H��_�2M��:�!�.Cq��CU� ����Y��LN��&I�>��_ܩNɱXΞ�=L"�p�*O�)�ļ��\�W��&�2��b�Qt;�Г�RR��֜Ȯ2.�)ȈqzĘ�?w��pU��,p��!�۽�!��Sd�0w��-Um��O������O�>HK�;�-�P�5S�F�� @mKܯ��a�:�E(��ۃs3�-�e El��\��]�L�n�X~���~�4:��sE���(H��&[̼�����~�r���1]]u�g\;8��q��PҒ����R^���Pe���cɽ��6�;��h����!�������W����l�0M�I��,˾���+"b�3�烶y*����RO�µ��K{ ��?wF>��e������D�g�v�vY�GH�5�ϼ0�rb�TT��_��X��4 �]l}��K�Q�A�Pmm�<%y@����v��f��M�ZCmә��\Z�p�����ũ��b�pRQ�Jtj}���c�!���垣5��,�y8`�E���t�.R7�]oZZZs��aҡWO��|���Sr:�$v�����c��]�핲dkHɰ~)�	ȄɆi�Q���0�z��Y�A��T�P�!
���)u���� ��O�^���ӵE�#�64`�{���#�Nv�Gٱ�_�b���G-/�P��kav%pQ
>E-�~ν��,[��� ��J��1� �����i��m��s%�z��̗|�P�'ֵ����c���굧�"��Y�?�?��N
��G���{PR�8��I7\��F�:�Z�G�t�چ���n�IYӀ�������`��!�sS�o����7���(����T�P�\���Gm�L}�=`t�٭r�~��X[g���_����AO#b��ȩ�"�]�������;��,�s^��>I�-�$��A~����z�Cy�:h+�H�;�}-wЋ��+�<�34����>��bt�,�C��8�6����=�h��WJ/�M�����-W%@m��/���vЖc|��>�d�$ :|���ʧz�YR�fR�lmv�R�7���jq��������
7����?\���i	��V���uv���P�����F [y[c'!�W���^��l����*�pO����;
}�Lx�#h���k��.㔿���w��T�s�dUFX^�u��<󼌣x[��L�ʢ.���(����Ga��i����
#yV�K��+h�h��cĕ����ᤐ@c^|��h?�Nz���/��y�c���/q*��+������\��
UU1YT�ȶ��b�e�<��f�C��Zp���줤=�ʮ�IΒ-IQa�B]���g�_�eC�s��něB�&��o �HwK<���?��(9.|Xo�I��n�x�v��y*�)������BH�p쯣(AT����=㕫�eҀ�4W�~]���9zy�03��6�ނ����y_�R��z|	6'���e�O�K��.�@~�Q�^I�;��w��[ɘZ�Q^��n��/����,d�����F��8%��;c+"ԣA��:���۞_�H����<��hF�i	uvCq�977�ֲ�;~t������'��xt�l!��z�!� l@��/����c��~WH%,<�1K�oQ蜭u�X���_��Ci�CK�N��S<�WV��p�^��o�_`4�<�냰����R��y�M��w(���K���OD��?�oe]�k����E\8zϽ1�r���)2ˁS��2Y5
�x�p��T�%X^Y����Wa( �rO2�Ƽ�J�%L���X����̓��rLJ�TF��`�:�M��cR�ɵJe��hT���Z�R�Py�`��o"��:��b�I`���#1�=_t�}6���N��t�P���>�3�6Hg4���Hv.Lc��HjS�Hn��3|�MF/��lYLs*�T`�߮�
�S�Í���w�}f!F1� ���0�~��9<�2���rQ�J�=��F�Ì�^/ɷȁ���9z��櫂�=���e�N���:��9�����f��2wm.�I���bە��(���d�/
0���[l/���(d˙��2���NpEQq��j��&w*1)���◢�U:�=�BϘ�Zu��@j0X!�n#���R� N)Ж'�Ȱ���i�;x��Ե�gQMBVW�<؀�P�D �vC��o��(��:�v�?Ei
ʸ� �kd�'j�
�?�؃kB<��Ŏ���>���Ք��E�.߂ �=ƝLˢo��&���� �^�K�8��-����>ͯ��s2$�f(hC�}~q���ZC�y�j�����]XٙP���3�C̼�0k²�Y��.v��ZD�C9�C�K<e�gB�
jΔ��d�X��8��=r��H7��.{p�:��5$�+�\���;���Z$�!M
>�j=����\X��Tl�P��IW^��[�b|�*���Vਰ���D䶻{��ւ{,�����Oh;ڟ���C����w��z[�g�^�W�V+.������>��Έ��lr���oCW��:�
�s8��`��Mdҕ#����T8	����ce�o;���In�N�fH�$��� �{��WG-�o[���{Ԁ�;��<��P��x�!	ݤI�fs3�9Q��>�C��jk�`��	��Ѧ�����7-1�g�����i���(�<� �y� ���Q�`;%<�_΂�¸�z5{v=�~*���}�[�71I$�����V���.t�Wn��P�r�m�&��F_�f����詒����*�v��%����f��Q^\�.:�#"�+���#���������v�(6�գc7�G��K���V��$��(|2�#��È���Ÿ�!`x$U�!PB�YF�2S�H9��@X��,=���HBN�"y���:R픀zF�FG��k�~E�>[Y�GT-/�e��W��N4�H��+;���H		T���:t��U=N���pb�k �H�J����g�[j����*����&�̚��H\l�u��ki�{��Ȱi�r�Vww��C��ԅ[�q{���� �O��3;���ȩ�����c
�uReo(c	���6c>�� ������<�Z�#�BeP��[������F�4,7��֪�v֍H;0�����#��&⹟�s�_op�8rɅ����E�M�n��"�$����<=V�o���=|<�,�t����ξ,; �D\�� �C�8�+�Y|�d��4�q��NU�al��ǥYHt�*�y{��"����1�24�'�Y?�@��yS�h��C\��g�Ť���2'@\��щ��b�.�G�1���HKZ�	 �R�lI���}ޣ���BQ��u�����Pa;��_vO��|ܗ��«�B���ƨ~�E��#W�����j`;e	 I�)o�0TlΔͣ�Y���h��i����i�͚9c� �W�gS��uJcӷ��g��,�(�����,�$��S,.��]���ftE�Ȭ`U**���j�} �oP@�P\_��H�ⷋ~v�5c����y�\�E�>��_MN� ��(7f��y*�����$��)AT6/H�GvF�)ۈ��ϩ�p�������dM�pty���M�;x5�Nggo'~'��$������M���13����C�)"�n�z�T{��d8>?z\�z���fc%�:
�űC{]��Dpc5ǁ��@D-��X��k5�i�IG"�ao���&@�%Oݟa�^�k�?y,�����U]�┹h��!�#JK��,�x�"���Rp���%d�?��=*.!.8����1��U4;�y�;�4���!��s����_üC��q��O���Nٿ�
ЭЍ9�?��`lwm��'��:�FV0/���l�G�Q`Y��sV�_#u36�7���( j���Bo�fc�+"4�j�<EV�0|�-0
��Y��Z+�D��2">X)���0q�#��\&l��DΦ�8�Z��Ќ����3p�nW ʐ	�b����<� �t:X?�����8���
�}� �EY#��״_F\<Y������w3L�>(6�TOe����Y ���I�J ��,,~��%iF�[R���+����e�{�ȉo$>�-��X���ͮ#�V�s�/T_��k����D�k]��=�.���Z՞]�]�b4y��l��v��zB���ʲ���D����)�'�wr�2�e|aװ�!.��;��45{�UU0/P2�8Ķ(�ˍ�EX��/&o�f��#��l�-25��.	"�����4XQ$�͎V�YG����N�e��~,�������H��fs�,����X�.�<(�,����� ���Vnr��4@���o��nj�S���kӹ���v>$�3L��鯞b���]����2��_���<	/P���+���R�:���y-�m�´饢]�7��sAk�*����Q�����T8�{r�2��WŊ���A #G�371�� �"ęi+?B�X2��s���,Rn�_�Ǡ����'�������f
�j��8���e��<���K~t� ��q�H8;���U��)j��|@�gw��m��:'�m R
�-q%�8.�LD1�r�3R	�����t�k�s�	̺fb߬�׶2���}"����%�vɎ�#���6��̸���夽w�g��<�O\2�j��i����>G@V�檠῅����t�����N�pҮ�����1�b3K��5-]Xi&�+ƈ��! �x�}����,���:��8���S�fz1�t��:�e�V{d�����Զ�#U9���t�Ѷ�a��P>4�5�V)b��|���۸�Ϸ�O��q{�Z ���	�Ӝw>�' �Y֢�H��Yo�}�O|n��_̺r�ԬRug(�4��2%9q]���W�	�4��N�ogB�Ԭ�N�=����D<��X�xM�07�Ż\W��~<�{���J%\�k�.��s 9O��	�@�m�:�K'���ei�	�����磙;��ۺ��?-_]$>iK��9<�:F��0���8��W۰�)i�iHH�N��t_W��h�ì.U	�P�F���|�J��{����T룄���b�}��`����42ܩ��	�����Y�<�˯�;w�)�e}����5t	WX���!����R/���u�ę�z�m�[���9��,l��`����O?Xk+r[T4�4ѷ���+�9�O˽���a��Q�� |�A&/�lŝ�dҔ�EژT�)7��7��M���{�0#,?���OXR@�rÑ�W��wV�r������T)%J�I�t'�z��nW4p3��l|�Ӎ�5���9H�B�܈��H� ��^Ʈ7v{�C"�H��OЀ���[)��-Q�v��r�N'����M�s][����Xcuk11�!t�3'�DaI�3�� ���u����u�t���ʑ7M|쩉\ڛ.�+�==·�1c�}yy�}^�ğGU��r��S�2��J�Y��D�l�or��G�xR^�ش#�fK1{+�[��~ژ;���&��=�_��Ģ(�:� >��/�p0:*uLe7��� ��o������$�V��՜�s��"Ъ�m)��r�ʺ�����0� i��^b(-�hc�xǸѤ��K��Y|uRZǳ��#�h|�q@�Ҿ5����Zc��� ����,D�c��m�G3�n��4^ׇ"�E�Pz�e�n�)F(]���% ������u�n@�bH��WU���iǫ�B��+�����Z�Q��|fW�	"�I@ڔt� H�S���߹��)�}r�tF4���lTtʍ�32�iQD�Z��UU�oί��ٴ�@���@\x���Ԝ����H�b*�?Mu����D���4���Yʖ�+c������M��,�|}̖��
��/  �%��	����1�f���.m�{҅�8v~$�H���'Ⱉ��'�:7��բ����d{�nž@ɵoׯ�s~JE7�P����c������Q�R��.N�Ƶ�k����^_�#�ۃ�.Qz����ìF� Z�e�K����+qU�s�ލ�QC-��h4�*�> ��c>%$;��]�q��3p����.���\06D橧��@hH�U��QJ6eN��f�2;Al�͓�Ƥ�p�-�}Д�)U��U!����\tØ��}sz�.����2�ȴ�l H��8~�u�V��S���QA.��-Rӊ"�d7�_U���5p.�Zߝۼ����9�M,���u��Ԁ��ΒVv�4�g��Q���73(w�U���tT��_���i�c��A��j�զ�,b^����m�G���I���� ���$�$^)p��x97�t�89"f@�m�m��]��n����aq �x����n�'>�s�iS&;j�̽�k
?���WPt�W'hB��d��]�OQjz�nu���OFVs �^�^�͸�F�n�]���xK��W�!+���|;LS�h���y���7=O�D��I�28�a��J��<Y+����`�RK�l\���,�R`fXX��XUQ�����3��1��f��x|�@�-y�8�y��5|i�r&�1rIA��	�|]��.i&T��b�j�1X��省;/�h���mOT�3�o�$�~i��,i����H�^E��@��\�:L�!���v�NeD�B^��,�\7�\�����8�,��d�7�搪�� `	�S�U�v0 �+�n
����ۈ��\g�b��4��~E�r��t�m�E�c�5�2*�sP2<*��Q�򧕬�)���"Iy;�	��ڽt^��
�� �>.���4}ɅB�fθ�����a��R�~��zD_��ݶ�=(C@�����P��YK��W�~g=@΁������]����|qք�nⷭ3��	71���ކ|Ϛ�o�H��p�jrɻ8P�m���MA���E��-�a��%fi���t�x��n��ѿ��d-jzv;�ݤ�>�1s��o�r|��ľ/�Sq*��#rI��Wf����ـ7��M��$˳Cb$0�
N��m�.׀%o�!��d���3��k--F&���,t��ɹ}9���iXt��}�ʔ���[�o�i�x=�F�o��7�������j������=g+�R�W��u���|~�-bfe�ᒉW�Y:���+�x�D-�L~9(g��O·���;�`���V��3q?f�^��7)�(^�z�XĈ_�7�X�tYG���dZϳǓy �]��!�Yɵ������)�����O|?l��]1���(,©5=��2�`�g^'>mH���F4�_�Yr���m��Z��}5aZ�	����.��Uy��.�2̫�P�{~D����������9���)
K_��/��^E�x�������Fue��r��0S;?�j�������2C!
�����V�lq�d�í`�ݷ�s�`�����~h�����ҥ�\���=��
�Z��ң��B�J�E(}�� 9��iF4e �7LG�:�HX�9I�p7��b�
����-�7�I܋��}R�[+�Z~myߨE��DC�sI�$��A����		��ٖ(�nB��v@Ƞ���Y.��D(��,2���5���A� ��hW��&-�l��!ĵ�ߜ�'��e���W�N�뤴g��^������v�ٞ 	w���tA��#{�IY�뺇�<�X�"*+M�jĀ?����qv*���6�g!e��j&���أ��Q�I:'9.���ơ��
&�@̩)US��Z�	&N*��kB�Y���$f��!��ڞ˿�+�&M-Du���]�Ĵ����S��k��q�fT��b4��h�9ʔ��ky�-�r��i����F�:�[ 22���z*��{/���~��'ϐ�*����$�{�㧖?�Rf�UeCP"���F�axt�y.�u�嫕�����le��K�v%$zE��y�f\�7���"��ebÏ�V����ԝ~&���}]��a�h�1��m��O"4jn��[��ym61��S��5M�=��T�y���~{^+�Gr�gdw�K���������iy�03�qb��8O�O�E?�L�����~�F+�6�F�뽠�_R���xr�z<+���bhTu�/3��]z����Q �^L�7��nȲ����!��zG��X��LQ|�������Y��:�duc�����a��ΤդlJ�C�It�'�ٳ��ȴ+!�B�ߘ���**w��2���/Kt�	g��:yHV��=�O��Z�E˦�a��P�k��Q�`����F�(�6��c�l�dhA���,���bn:we������K8��u��v�P�t� C<P��RV��x�R�,K���#G�&��̜ꓺ�
��O��q	�Q3�>cf�8�(�	���z�.�{tc�%׵#�ξ�.�u�o�"�n?M����lfx��'.�c�����%�њ]<δ��fr��*-k
��ѡAkM4n�n��X�1�T�P̭{��D�l|��'m�'�[���k$��~� �i��=�(��D��Խ]<8����(`M0���ѵ�-0�L�.�2�%��j�f�S�x�hh-��߫|&p�;����ˆ	�O�B�(#���&����֍�#�0�M��v^@�� �Cr;S�Y��.tZ4�+˧�`\�2^P�Q8o`:�Y� �2�	��d���5�����9��`�1ĥJ��C�Kb���xg�'����9w"'8��Ak�C�|0�d����a=	$�:�!�ca�
'��}eK�h��Z��;���p�=�R�k�m�ȹ9��Y�����~��=�k)���L�����XU��BT3����_�H�[bEX�ك�;�������7�V<�53�B�o��l _�u���̓l���	'�o�&AC�4�[9d�M�/��,�\�el\��� �m~�&6�p@��jYq�O��!�������v?�YP�b�\���ۤ�Vwڻq�a���K�+�Zo��",�S^�-�VQ��f�;j?m�4���ZI%�l�)a��\�7$�zPO<t*O��b����m���ݒ�Nh���VT��F�M��P�d���f�*	Y�ٙ�y{�+�aH9*;�q���Eң|����%f����� �+�@�s��
���7�6��-�b��E�R���.����Wv��2���-jc:$!n�$@��u����2]�5�h.���6$��"ʿ�I@z'D�}海�xcŝ��8̼���,]����E�l&����s���&=�;;"���m�Id���C�o��6�M#˂�o�W����_X�J�９�G��ZFN1�jQ��d�w��5(��3�L���ww�MO4\��F��#�C�{oP̬��r��V�x��!)�}Q� �H��2B��"|��1��ڨ�<��($]��Bq}0��{�:�.C�H/͌Ӝ���v�� �bx6�����*Y�t�P��<��\ '3�T,��$~o	�b@U����&��:c"짺b��=k��>zd8u�8���"��x�KoqƵ ���jۯ�/!1ŨÙl���/t0c�4D/@	��@��D�y(J�d˲\������P?ip����l���hTԄ��.����R�]嬂���>	X���p5J��t1{�� ���S�q�`�Y����9��['^
�H�w�(P�����z1C��rG��2l���*�������x���h$����ô��򸚒ҶR۫������^��1���g�t���tf���deA�X0A ����ӖG����30�6��E"��jw*n�Lt��B(�+�&�}3S�43Q�J�|_��,���c�G�9i[/%D���(�Wqi��CuH4:³�Xzޙ�i�6��K��TZ<' �,���
if�8oX3�{�",�_�IWu\�����^|�� )�TYI�I1_0��0�s�vW��&Cu��h��=��h|�'�~pT슡Nȹȕ���}���+ʘ�h�H����u�{f��+�Y���K���;9��|��P	'�iX^}��}[���CӺ�<����I��K*�a�`�nǷ[�iT���u��A��"Pͧ#A�?}��s��8�ݕTRkc'����S$�' �u	�֯ߴ��a�j0�kߺ�U�w̃��p�o_�A�75#
I�<�YoW����ӧ.	<P����ɔ����y�߂�p���è������'ϝ����D��s��r�����mi��hΩ��5j���`��3p��S�a��d4���J�&��l0|��xc*�����
d6Gt
V��v���Ŝ޷_7�	������[�p�c�;��/�z�2/xw=>^��owİ��_���=�c��U��	��ޛ�X���r��Lw���S#ru1780�b���T֧s�d�pӤ-v�bfɋ��жU2	�M�� ��ƨpW�r&Y����<�SAJZ�W���٣��Â���,L(�݋�5�{pP(����噞��Dt�c�k��Y%�#�F5���P�;��l�7';b긩W�5*v��'=�Z-��㞶< ����p�JS��I(�A�_�)x`�E�J�oQa�l%��$�Ǯx�l|C�vٸ���2�(7݁�9|�?ޏ%��r����21`b�!	��T)���;���s���P�MS�HIcbs�����i�L|��G�d�Y�yo�j#F��N�%�=s���lM�A9�1 +��Kٗ��l���@�l��V��S��OM��T�ز�h�	���m- i,3�u�� �ލ�haK7�=�xDuP�PcDI� F�|�}|�:��� �C`��\]C1I��݉��f2_ʱ���J��(���d��=��a��a�ȍd[�/S��'ٳ
,m����]���� v��T�zA�$���r��@���V_a^MEM)lf�a��w�*��(�:{�Z���0�t>9�E~��%^��%=Z͒j3�h�
����[7�D�I�"�,LdYI�b����"ׅ�z������H�r�f��$����A���-$J� ��v�Aa�bӼ9;H]�Z�uM�u�]��B�����:��,m�AW�*<�Z��e�����A�~�D� �`p�D��Q�}�����B��7�	<�U0�.���Aa�8�7�r# �z���b-�`���4��Ll�����1K(�Cu&�5�ə��R��}���5�^���/2��+�m��3T�����+`���X����RSJƞҢa�G�7?�g@&�/>��^�|��{�[DD�A��0�\��+9a%u�՝�S�<�/of��gw%H3�9�3!��ԍ�h��l
*��͆�	�P-Z��r�f��?OI��y���-���������>��嗃֓1ݓL�G2'7�ͬL�o�����՘���4�UQ���An=ᾞ��22�߀���&�@�$�~�6��{�uf���ˇ�5���9��nV�,4���j���M@_?
xQ��!�gQK���3X7h�apz�|�n�^��Bbvw�).�Ğ\�\X�Bf��Y�*eR��w����PY�;Om�~�~r�Q��-��@x��/�лҕ�'�͞�����]� s��T$>�FC����^�c'���ڞ?l����@��:<�ݐ�]x�T����i?A>x��[f^�+�F�)��ߛ�|�x"���tiv�l-4a n?����3�8W�>��Fv!W�hH�T��/o"�������B<�u.ɸ���P֨� ]�JI\TQ컦�r�����fql� �*N����0ڪ�qt�rfk@p%���ΨK�Z_TǧCF�)��h@?�#�ҹ��.l'��%Iv#�)�!�g��37,t�����,^�[Cf.�6���%�n�dFp������>��ZOC��	��+~���E���P\ H�o�Aee=|$YY�y��}K�v�����5P���|������mUׁ�(&G��O\)g~��h�����S:3�����%�W� 1E��N�A5�t� �tx��3��	͜p��'l����yx�_�1���O믇�ߠ-�.�Q�_հ��ڀ�<�7��`�,����+,D�q� �=��+pVZml�4���e��~�a���¶��"=�.�u7����K����լ��د�C�}�Nw0\�GW;-�!|uQ�'G|�4#���K����;+���7'���^٫�T�F�9R$rRUY�M�͇�F���n�%-&�+ע6	sޕe�[�镇�=-$��Ԅ��gM<$?L|�N@��fz��`� ��z(<J��F��u͗D��ӑIU��D!O��p3�e�f���ٕ�O�i�/�qK��������_��6sr(�&N��\��e��P�5fQ͎�S���ќ����Q�pk>��Ȧ" ��u���Z_)�/�)Z����.�����jT���(�vp�x���0(�Is@�i~��4��Q�s�A5�������#��]p���t"3u#���[���B%4���TTM.�%dE'�jcM��IB�|�CsC����x���ֹ�?,_���݀��ߧp/ 2�Y�;4c�����<�䴅j*s��h����
�䳍��Q.N{�
Df� wΨ���EC9Ѻ���i^��{f�[|��3�7p���� Ij���x������$�*�>��=�x��,��Dܼ�Q}���1QL�\t[�E�@H�+]3��k�Ui��5u�ƉF�B܆�d��?�m)���ʊb%�l1Mǧġ<����uE���O9�=�q�6O #Q���� �1��ꊖ/��FN+�%��|���ͨ� �'�xgF��wv0�rz��ڤ|�Ei*�kd�z�zv�#1έC�������?������P�z�#\ʻ.�71y*�˾���)�9Ly�/"i�62+p��������_T�[L�<����&�#���1�E6Ļ��R��6dT�^�ߡ�}}�Y�����bW��k�}#��u�=�:_����b��k���^�][�={��G+��&� -�@|��9�����R��e�J���g33�B�:$5���9���3�c�.�PڄR�	o�}���PP���/Iq�~*��1ǥj�1�~�jY帩�C�rX��?fóF�����ٲ��7Mčx������4#]�rM��N��$Gb4���}I�SY��Ӕx'*{�e�s�9E���ģ���5���]Y>���i����4�F#r=�H�̃v!����~�}b�(;M���j}>.�FM���y���P���m��wB�Z�N�Y��l��Xox�5)�l.�p�&U�f�N~�ӑ��}l�e��8�߁T�w���������c�U�)����Q�{-|65�m��p��8!_I1BS�&��%���%4���|T���"�g0b�g(#^����hJ�9�����[՗h�X�ߦ�tr�@S�бB.#�Q�,ˬ�}���*��ހ�^�<�tx�`���e�0�9����58�떚ۺ��$�Cf��hwbB^i����F��u=c�	i=����+��:y����wdg8��j�Th��|�kP	o�A��d5o�x���t�((�U�	Vw@��E\�`>%�o!�8�&���[��2N:��2:�C)��!t�Lߖv<�St��`���D�� ��-Ծm��j����=78�2ʍʇ<��.�ҵ�u����s���	��������`��62P��ц#g�W0�|d��T���9xZY���ÊX��Z}Or7ʒ5+� o���%���}��+<�ˈ��^�͝�V5��� ݟ����E��0��V˩�i�oL��<�:b7�%а���A�Ǚ����&�.�;�p�G�9`�R�'<��Y����	���mn��X�{�O����lq�$) 1�G!���Ix�Fn����~c2f�]��(E�>]��g��V�Bt���"���G)J�)yj��qp�k����c�G��;Ú�A|��]h����m��eA��[����f�Zi֫�
q�V<�>��p�$r��<q����MYF:k�z�u�2~2������-����d^O=R�t��\�]�sEc����~��>Q�?א��KRٷ�O���>�C���!�����f�8�3,=S��ӷ�x^?���O��
[Xz��1��)4۟�md�u��u�K�����1�I��\��A:y���Οҕdr�v�7���m�)AG)YN5^���2C��i����	�4���|�9tI������8s"��}�A�<�I_1��^$T����ޯ�M��b�(`
9<l���A5wq�UN�>D����F� �^FB��J;���5X�{j��xW�_+����m�������*�"�_4=Q��TB���"�*�ز6�r�E��J�Q�׭��cv숵m�t�1r?�%�i�z˳��X�W��1$6W��G�[�
w�_
�楲Q�snaq����W����E�&�
q���wwMd�W�gn,}TWz���$'$^���;2���ۏϰr�����F�,g��s\_����[�7��s���f�o)�1�4t�$*�gǘ�}�L���RX����]��������8��ܧQ�+}2�2�t`$��n�_�_̛R���yL\2��tiY�N��yh�sۨ�8�Ը�]p�g���6v.�i[�t�������l,��D�
��}���ӛ��#ew$y1��;-f��WJ@N��i7��}4/��(�(����I4M�"����k�y�Dh��������]�%˭^�#��a�ZD�"�olvN�OPkD����<��<�3
U�λ�����Uv�KM��y͎�IoS�M��E0��� T��q;���7��h��[�3����>��g�w��T��I��l��dd��8!����ם��~�H�x&��Bʍ@�x0�R@�׮�m����N�K����^���啸t�2�΋��t���ս<餉���!k2���\N�qB��{��`[��P�,_d)!��H��Ӂiwt��G��L��ª诓��T|���ؒ�3I�2xW��B��� {�Y�,O�_6/|��qV�^&�[�aL�����i�yF�x�Y\��cORQ���h-� ���R+�<����{֬��?*�Ҿ4�J[a��;0���FFG��{�}�v�	�+�7"a˺���x"e������Ry�%A���3C>���܌��Q��%I���DF����2�!(	,'�|���<e��v�C��^���P#�_� ���X�q���r5~⫺>�Uga�v���5M�pe�V/���%��ظ�����ƹq�A��W�@T:�/%0_m��$������@�y���}hq���N	��\2���ނڭ���l/W0�(8�%l:�?�F����X��*�$z������%5�������������N����UXf/�Q���H�G/����JV&�F�g��Q�~�����ex�>�ܥ���2�q��q��	!aPD��8�!�n�Sk�<�fEE�8���=��D�ݘ��*3�+���-��yH����c��w��z+*��������e�y�������1�tI.��U�-���y�8s��"�'M��bxe���\zoE_O�g����"0F��+��P1Y�I��!�O�¢�g��to�j����{x�'�uR�|��g�X��I�;���!���O����[17e�/(���H�ٻ�ТöE(��+����Y�Դ���/tL�u���i�G��3�7^�&�w�㢖���+v!3�C/w޳N��D��Y�<x&��e�X��
 �n&#dL'7�6ǈ6��Dd[�B��T����ǉ��ė6�J�����Rw-�b�.hҼ��D�j#��ԇ�,%B�q�=ʴ �<c̭0U������`�m�e�f� b��_R�e���ĸ=�&�M�%$���	��r���6�ic�_��5�L��
yv?	��vN{ٞs�a_�ZZѳ9���]�];�+��`Z�_�i����;�0�S�� �}���*�Vеz�"���b�Zn^VV}RK>+xfҵE�s���0�C9�N���h2��ȡ\��O��v�دt�n9�t��9x������/���K����5��3��{&���
;�bK��P2�M�LZ#�X�kS�y���耺�@E���e���&V�2� e��,)E����@z}Ϩ�����m�obI�{�*m����d���Ǎ�c��+?0d69�'>��R׍���-Z�fimXٲ*�	j@�u����h?eޘ���{�X��w�If��۟ ��Ď�w:����t���`9�i����.��8��*$mbʇ���8Z�T�Q'p���B��'���J�4`�����M��4;�o��Ӷ��S�~����`�9~��a�[��t�?X7?r4�X�hA�;y�r�SOEN�\D��3��c=|���	H��?(wĻEg��u�j�PQ�:P�i�nJb��X՟B ��K]q�g�g�qα���{�	J4��Yu��+���)"�� D	�kh����_�M�m�{�>ʓ *4�S�f3�M�#6��_�����iH|w�ۓ�O��@�2�!s*ECU1��{��b�p�)^��F���}^�D�]b�{�kǸe��a�����n��:�� تU	�����R�u/���!,�ND �7�����E��"K���f��GZr���ْ�m���������ejG�1 +������[oÚ�Ck�0�Ӡ�)��)���V�\��|����w��Ƒ(��ކ�t+�)��z�r?��=�P���2td7BG�Au~'�n ��E�ųe�>m�pE�V�N�~�s�����6V �/˶ @72$���Pɰ��I�z���f��n�?���!�HH�yXVEE�J�/]���	���L:��\�#D/=Ι��r~��s�V��49ʄ��Sv���oR�Y������3Nz!�u�1\��9��J��ӡ�uB�&�]!�����A�ؕ/U��<�dG�<_&�k�a���H��W����k�/�/qU��T��H_5���E�+�H�U�0=���[��Ѧp�f)���V݊���K��ox�ʭP˱黠�J4kڏ���Y}��]����2ݞ�F`�I�M�Bq�����\r�{_7�]�u��x޺�}�[�q���p�E���B/����ׇ�ຆ�^�p���,<��k.^�f���8�F�ٵ�$��]�b�8���Mk�`��i����O<廆e{�����$yr���6
857%u��cL���&��J��ӳ2'�.F8����b��"lCxE��׭���#Xu�A:�y� r2oF�<r��<?�����|���������G�>�bUs����)'e�9n�)�)�ق��㧠�[m�)$e�E���Y6��n�r
YP��P+��� 8ǵN��'V��=4��W�C��rI���u)y������!�md��j�N���X׾q+w<{xp�$��h+�[нH����)���Xٞ�;����&k��BM.,�[� mEA��LYg�圎NL,�(~"�T��GF3�I�?�T�#�!\2֮!�%M�+�Zq� �V���Hk{����fr�j8&`�e,��jd�}~Aèy�"Í���=�3��R�l���HV�8�J M��A0�S���uE���h��c����6c�w�y/9$��I��d8_�0Q��) cȷ���V�d6�.��kJ�f+ q�ܥ���������0"94Y�M'J�h��ƴ�ѧ�Ԉ2C8�su�D�1�Q�Ǽ:�2v� �6ߋ mn9m�s������� -��U�Պ�#r,NxS����@ &ѧ�:^�g.�I��ة_w���E����{��?ݢ��[Ӫd���	���O��d&7��s'?��5p��o�h���(5]�8�ٚ�<�Jʴ�WZ��~e��K#��#��1���\h�[7�j
��W	3㿽�(�iG���r�2V�@�#K�q��w�ժ>��dti���%&�0+�2��6F̣�����G��i�'7;^��@�&�v�Z�G���vצ�~��٠ju�X\���O�C�H�ă�w��ڬ58����Խ{p���O��`[%|���pN�h����S9�·�䵾L�,�"��t |����O���uO0m�<����#V�Q���t)n�7GׁA*��c�����Bz�8�����?ck���Vy�()�0��� �V݄&�%�{�c|��"�x��J�Y��H;��ꨳ	|/�7��Z����N�J.�f��]S�&�(vX��ZU�0�s��"���D���t�WuG������b׈U����2�פ)`������g����W�]��k:����UZ,�:\�)�$U*J���D�..n������g�}8��>����Ҝ����!O����U!�W�&�:��n�Wi2��픖д/$Z
��/  �O�Ki�o�	(%�(�áS���R�?�$��1W���2Zpȏȁ��,ɒ�3a��p���VD�q
�g,��NX�mpS����.z���rT���Č�l,�J1�"\ʾwj��'�aV��5��g�y�װ}��1�y������ŌФ��δ_��ߩ�b���h4�*�> ��c>%$;��]�q��3p����.���\06D橧��@hH�U��QJ6eN��f�2;Al�͓�Ƥ�p�-�}Д�)U��U!����\tØ��}sz�.����2�ȴ�l H��8~�u�V��S���QA.��-Rӊ"�d7�_U���5`'w�}G��&������*��ʟ;a4�_}�>K���� ��9�$� ^��1��w#��Fu[d��9Fmx�u�<W�=��7��E�.岍�+<��@X�)��^X[2�H�����8҇�f�7S�w�Ց<��n	,H�a��biu͞�)e�YE\DŔ^K��KV��@y�������t��vx`d����oK�^y�Kf�޶L0��y��@0AȞU~�;����Q�"��ͨMq�H?/���Q�7����x�}���p 61#����B�`X��b����\��!��ϊ{5�]��>tc��	15p[#�ό��I2��L[%z��Yu���@���&܎�a� YtDh�"��r�S����V�c'�¨�;�Y�0l]�.�!Y�o���n�~/d��`X���^j#�?ьI->Y,^�$�2�'�V-@�҉���>�m;4�T�7z�J^�V+̬��:�z�jƃ���f��asU%��[�d%��T~C�k�>70x�z���J^J�X��h���ۑ"?M*o|bu��
�@�U��T�P��Q���3)���⤥��n�l]
�� �n:�M<m�����]�wǒ�+?^`��W��j��TLB��Н�.5�,)J�;G9 ���#�)���8�g��3�-[`������&�3��)IL��`7���.mT98��FD��o�Z�@:�傓rx����-*�l�'�Z�*��u��*�,�+�p�J�&T:�6aI�u}c��q{fl�XX�1li��v�{�G�30�H�U������Y�;=[B��)���|C�A,��O��@g��C����v51�x 6�L�@����VJi�(H��}̺%b�TAg��|���TZ[���������*�i׵��9(��� ���k�w5��S�Dϝg��+1�͕&���\1/�dg+i��b�ӿ���.w_;�q��M�Wt���JyI�<v�_.g����0���Uf5X�M<!Z��A�@] 0'��sp:h9��Rc�;m�4��/�Ԅ~*?��ߪY6�I�z	K���2�i���5�4>D����|�K��I�g��u���\����|ђh��:4	�
����e�i!T:C^�$��	���� ݺ��͠���x��DՉX@S���Y�ԍ��C���/��U�B�P�����]⌇@g1�+��z���|<��=���a�ք>��.bf������j�����͈�KF��@6F���v��܏�*N�X`��dh�w�4z({��c�`���(�%o�`/�SH]���Q��X���18!����G����st��{��� ��)c0_��A�n���F�xR��)C��(c�`���=��|�ܭ�܉N�p~�&���Jq�����\���Mj�&����DED��ȥg��pח¶+a�k������z�ղ~	�)�w���S�	��$M���{؉���W�������MzBW�m�����E�(@>x*���)+�����?)=w���YQ������f���������D��L�{���x)�A�r1_@�`(ϗ��b/�Y�-C���D
��W�m�y��δ�m[�=�,��<����P����P&�3���u:�ZA�N'�i[�%]�=J���Ha���*����Zժw�#�G0$T&����k���]5;�%|�6b_�"����l�)�M{����D��N�j�#1��g��|�~�����8BE�G]�����]�cQ��%�d&>7(X)s�^kZ~\,�}'���5f�c�ZjK9H�:��$��6��u`�b�o�l��+��wH��d[k�#)���]`��6�r�VK ��nH��;	��N*3����	SR>KZF��^R��<��>oOFl;�9����P��ӣ�Jي���7�� F�� ��qn��ɁsS��� �j��<$<�Oey>�d)kyNZLJ��F��G�?X��$?|��d�S�z��f���'��8��s���Ϗ]�K`��LD3���8�K,�Q` G��ZV-Fj����~�/p~���G�t`��:b'[%���m�Ҋ��G���2(�L�k9ৈQ���suw8�vYL��]�XI��#�2MT���Lm~��:�x���v�ٿ����_�~[�E�V��<H�tOP_����Q��7hۙ���gJ�J��B{�2��S!�v�21�KfH�0�Lo��)*�~�(ϟ�D,t$���㚫��{�㊻�)��Bj�r^��}1��NA�w���~���ʷ�'~���z0����u��!x)p_�{��jF[8��w�YT߉s�a�,�wٴ���Ǽ���g�����/G�TT��f���s(IG�{�b� ����eB�p6^����c3/�@AR��f���a�*n��`�e�<���eH���}-�w,����G �eAJ k8Tw-iz(��� F���a����Ӄ�����֖B�G�}��y��X������d���-��0�N���dql<���yV������:��$aeR�4��������ټQՐ�R���J}u��'>B}9��B���-�l������tz,Y�g�e�Oe����8�	�N��{]���Bq.�v��z���֙���� �Ƴ+u^*��/�b�k��QmM�Wc�+�8Z
[/qEh��1�C_��zy��Nz�!;��i������2�O�c��k�f(�����x �<�bz�+��p����v8�a��h�vlS�;����q���CStyȜM�y�L\�&L�{����i�F�|R9�I>rR��sܘ��d��1���#$O�B��/�`s���m�y+'72G:��u�6��Z\��<Ocy;���v8��|:��	;ӻ��5X�����o�Fݪ�S�&Y���uJW�*�������R �0�6�~ߠrP^Y�W{��1��~ 0��ͤ+����!��v?����1'j�BT4c"�|����s��w�BH����L�����؀�7ڍ�ڔT�)�ӑ����M�3U���)K�����;T[��k}����F���"/J7��1��)LXkg�@�1���h��z��l6J���66g|��(�'�k^���>aH��w��֢��2����\$w�5� ��^���g��y�5u���e�̶뻐���6_�D���儾~�Q)���}D{HT丸�?�Lh�[�n+���`lz[��.�K�/�T�����L��t����YK{� T�WK"��V_h	ȡ�^k��`u�ן>$َ��	ߟ�l\=y��	�N��
�k%��
�%��
�¬��t������/<)���2��g��l֚�>�F��D�l(���ab�/�F���dT7���%�^ ��jffx�m�x��.n��#���:�%�a0��,!��\l ��[����@�f��g�N%�H���^����e���"�Js�Zz����?5��C,��4�Aٸ2B���2����h`���]��������_�}���YTQT|`@�sq#���P���8�UR�[� ��jŠ�9����+�0��`p�U�r �՘s�O�17�d�����/W�{s���_�����8�E�D�B�' B�8��� /TB��ƣ�W*��f�~l�GW�$�5�c[%�]��U����������*��ͦnO��P	��E�%����Qb7���1��ki8��� ��	��TCo��h�Z�j�4g��ګV�������ǣC�X���l���ǚK��̃���Y��C@����??5��!]u�4�~�t���Է��Q��VB�ȻT�U�0�ES&S��2�.�����}�oM-Qhk�-5Rz����T����!e��{�c~�~Wz�y��đ�|��Ζ���s���
�ִ��*�".uQ���f�A�q�B�h���q<\��/�x����{$)�N�a�)B۰�k���
�=��V�m/n�����׋�-1�z,�m�M"�\u����I(������F4`��űJH�jC�@�-�wˬ�)0�>��Ұ���������H�u�t��~1AM3H��z?�3�Z=���)q��q8o� �Ei/�`�;Y�K��Ь)������|@��@�v��թ IɆ˦����Y�����}G)��\��įM� �Y�Pj�-U�h�����F~0?,��e�S�(�[�qUA��&���N��MS�Aӄ+G*�Uj�Y�$\������v�g�7�Ѭ��!��*�t���G_4)�eMK�������%!ᣮSXu��H~��t[������U����C�����)�@�u�0����G�dg3^`�����������X,Z�%��T�5R��S0�u���W��)� �R�Ɔ��gj�>�)��)�d�$��Z[�mAhw�>D�������c��>Vs;m},T-岮�`�l��@D�����I�YO��UU.��/^
�$��0�F.��49ɕ���(&�U{
���nwoAǍ4���.��y!($�uI�r�T��/�L����Ɓ|��|*Be4�4a�~;W	��
���i��L�!�v�P媿���o�J�if�����KR솉��ZI�%%X��B
k�vOq�YN�!�
e�s#wC��k��#�*vM8����W.?�&��=��Bn���DA򡔂I$U(<�  �����I��ˠ�'��~Q�-�U;�(Z.��xڏz���YZ�*�S$�g�������t~ւ�Y>DQ�ŭ��?��.�OY�×�sn\ D���1������K�nۯ�,������ŵSEf!�W�d�W�����<s�ܾ���M����Y�M55�-�a�|l�L!p&���*Q�,���˼��*&��j�"�ig:ԁ3퓝��L=&Z��^$��Zh���O��9�?��e�a9Q����.����Ò;o@;��������Lc|�m�V�D�MJߖ�L�4���|+%qRY��M��FI�2|����b�C��;��Q��>���'��#�N����u1���{QF�_�p�q�5�+��5����ۿ�RN��:�J����q�$��∾�5z��S��P�0S' 2^����#�Ǵ���>����F���0ţ�.�(:P|�aK�lx�]}�����^j&zI�p�,@�+{⼀�7��	|�;lVxh���(�BQ�����gz8��zF`^��=en�y����>�K���>P�����Q����xO�8�Q�bO�U`���k;%�&h)	!��>{~��ڻz�`jaS��	q�ٙj��[��e�\�6�������*~�7��P�e)���T�;}�X>��}��ʽ��Hd�TP�J�H�o���Zt���;Je杙�q6�O�AW���\vb��Wb�L��m|R�zm)e�y���[|-�[-|o/S~5��	+N������D8�.�u6q���Xy�Q7'Η�#>�����{��+�+��ͬ�{�D.z�k`HZh���mϬ�/�F�b�b����hg�
Ľ�����8~�[����#��Z���Z�_<U&Ι�U��5Fq�&���7P�{�5��`�P��,���NDFb�` Qʀ�'h6.�Bdx��+���p?�-���Y���Yl�)!�4��� 1�|�͌E�y�����~R��#��-�1��`g�F�P�m�㭽Cq��xZ0��i����o�p�ĸ؋U:�K&�SjZ�#�c�F�H��5+�(T�R��3�K��a�r�p�����q\b�\�eDL�sYR����d��K�@�iܠ��P�I2�[���s��E�h]s6��Ql�xl��~ؔ%lY�����'���Z�z�y@�h�/��&��y|����֚�8��U>hˤ�,�a�7O�f����{����>z�ë�Q��,�U}����T]�݆M�z]�d(� ~:�G�͔V6�⠺&�������o��i���x��0�d�����&$;�6��1۠$�]H�&���Gz7��܄��fk�XW4��������%��Wʉ?�	�����'(Z���"���\����;	-T)kB�ݓ�E~T�<�q�\���3�6��	����$g;�/?t��^Q�%!�i�]���@G����`�?rw�#?DH�C�_.��Gj^����41L�Xf$^��m����m�|�;B��Ȏj���=/|$j`zp��=U@t-p����H��n_u��_Y:��Z�i�y�Sv��6捅�,��VI���E���f)��!`z����o '���"-���t�n]��(	����]��Ն���А��v���`D��Vpv_�A���J%F�q?��/����(Qصu�$���,~�i�jA�e����7��G @#!�o���r*+�M}��j�0�5��ۋ�絠nk�:�D��'S�$]*;����ٻJg�9'UU"�114%�0�!<X��Ԏ ������7O�����<��i��	�O��k|?�m|9J�mQx+}���zrm���.�����V�ML���'�r�ǫaȂ>n��mߐ08w��V�>�b��ǭ�	�w�u�q5���#?�k�Ϭ@�1±��G��?���)q��v�}f+�]��5og�I{��󿴼��Z�qi0d�p�Oή�x�Z�$S�=Lj"*��u�)n ��"B$).�������A�G���w���s�ڧ�Պ���sc�dg���8f�־�HA�蔛D���P�O��Ɖ���ƜB���H_;:#5���
�*�s)���:W^f�kT�(y�J(,�8Ʉ��ǆ/Tݱ�!��q�=�C��#,y��i�YX�t��O���#v���@^�k~[)�[o�%]�čjAɰ���5ozF�=��n�Wl�z������8���;�zNw2��ߥle��\S�ڰ�-ͳ{e��3j��\�`0be�����`��;xc�֑�3�;�R�2�+�;��m�D�j1&>	�S�S���M��3Q�ƀ�O�;y��� @JB��df�JՠU��Cy�����E�Jݸx�>ٗ/++�`>�8�d�d8.�B�Ȩ!��e��R=��	�Jzc� �zF�x�n��8$s�uDmf��9�O&����J�n�{����7���Öf��]��1�4�f��.&���d_�����MvR���ו��.��['��κ�<vG��2l�74�����>2�wT(��Ջ[�qy/��Ǖ"�s �!	2|cҀ�oǾC}�~���B1��P��5p�y�
��Hq��I #��:y�r硩�샥"�����yƇ�g�����dE%dl���J��a��J�5��ҺL�0	�G�s��L�.���'��!�'9. �݆!?S�/�R�׊�@�H?Y��>N�_�{�bTLA �[�#�*�[�`�Mh���!����t�7	|M*S`�-;�����Oz!�F����bb����]>@5��g�*�V���N����N#J6�{�m7����Ņ.����$'VL� u��]� 1 ����0����rȄ�ُ�_2h��31�~���?qa� ��ƻ�e��L~F8�|��E(�m[�)JV1�x��
籭Xjs�S�q
l�[�rU���ѧ���C�!�{~3P��>�������&N䤰/t��R�@<���o�s�E��9��r���l�mD��t��f��W�6+I�Z��:�Ŷ20Ww�5%z:Lq��N�a���fm�����/�jy���:3�i�OE4�P �J�:5E�qB��7��)��B���|�y�o���9�Q���p��ʡ�M��GpL��	lz�ngS<�N��_Uʮ��~(n��ӹ��*�J������'އ@���?�݂M�-���?~�|�S�䫶~b~��s)0�W�8Zy�[�*h�'JuG#p�+�v�B(��"��d;��� sA*�j췆=�}�@q��x�͍�0�#�|X�MX�f�S%_�5v�u��p�'\�yk���W�phl�~��mu.	hM_=ǝ�ӑ?/9��[��q9��]�٬��@u�ݨ2��ގA���~&�SF�'��.���P�W׎����#�'� ѭ��KG�t��]��~l���j��۴�AQAIQ������I�Y��ҿV�"܂�w��+yW����<p�DfdI�!�g���b�H��s;q��ݻ�� �7��=�Mܤ�[װ�R�秞"�s��;��Jgע@�MQ^���)D��e5�g�'�W���z���!��5���LU(��@�d�n�	�/���W޵�yO��%v:�GSE0�}���ڀ�#r����]i`�9`)ݩ�G���dQ֪�w�K�`��7�V�M2⏍���c����h`<�^z?M1�JZ}&g��Q)� �-[������s��RC)�`��AS�[�i�{�ߕ��6�������g3ƭR'�\{��m`��L��;9�=$��#X��R�^�1�o��N,U����?,���}�=2) L�ｧJF�<�f���yN ��s�>U���Ӕ�~�f�c��1�X�а:��>��χ���R}=.�}��3	.P6�c�6)^�WIAk�y���v��D�fAz����y 
:9A2hq X)�����=��|2���Y�D'�z�m��B�<�.�/�.�2RV<��PR�����UɎl˄탶�@��Zm��m�O���H���8)S�,��]5j{!f��T>c��[p�s����5���2�����w�%V3W�;ILF��=����:�T����Q$���������E��3����6d�a��)����m�~k��P�(L�>^ܼ�)iKmzP���h�'�������6I7?�pg�r�:�a��D�]��*�,�]њ�(���M�C�s��B�	o��:x7�0���M��]��jM�$�TP���@@�@���eEFq3L��:��q3=�F���g&$��^���cJ�[d�tb� ���]%8]tl1�n�"�z��'�#OƼ��|�e�)��M�V��e8�`�����rf�%�嘃/��w�ǟ���H��=���68�\��V������s�m��CԹ[�5;B4���$�@j�ddl��,��;;so3�h�����)�q;h�j��X���Ŏ8��A��;ec��s�⮩P��>�w����Բ�.�z�	�C�eJDr��^��ܜzu���|����l��C�<0��nM<5�{%���/��$�պ�HA�O��5rԦI��f\��<X���U�H��Ϟ��{�&����=��b�O-:󬉁F�Ш��ѲX��H��8�ęG�8ECځn��C�A�r?�.Dn.�ڞ���"-�ϰ�b�c�6H��Iꀈ���`�ixሑ;PG�����./�ʎ�8���6A|���w��G�W�!,���5��%\b����
nC�l@UL����|+��ѡ�S.6J�4l�u�5��·-����W�SNG�苃͐��,ٰ���ի'M#�z�y&}\��0T��͝�^��9�Һ�T��Z^�,��6�oJDb_�Ö[ޗnND�lgc��e)���;�SՓH=N�+�a�x��M`�n�3ٜ��yڽ��P�����a���4��*m�͐*�Fe���#�v㠔ޙ0�!?��+��a���l�~��:EXQ���R��a'�� a��*�֪5�͍|��ƻ|���M�d�De�g�rA�>�-�>r���M9����F�������4Id��
9��{�TD��Rc-�Λ
�A�h�x���^�r3X�`�Ƣ��6���sa��0bbq��.x�#y��v'���S�Bk��=Wܫ�y��ծ�m��}�1�۶�c�E��e�C[��zAD��=��A���R���]�k�\R��{<֒J�/���.B;U�Jҹ�S��1��l��0��Hœ�<O5�����aLIC�+��ټ�?Zh4_B�	�*Iy�$ƵjMh��?v �ȉk?���X�G�i�.ܸ�ţ��&�Ѣ<�(h.1�E
%��:�ɗ5!�y� W�tT��Y��`w�Si(��g��l��ҩ0��qg�	�I8zʘ��'+�!z��9H��2�����c@���8T���<�����j��
��Y̿	�=��\����YcN���;��	��:h{��P�k��J;�Vӝ�o��h��|IBv��[��6�g��)��`�"9[g��"��R�:^[�[K�I^p�Rr咂�KtL��c�[�?R�����Jy9����X9�jO�6�Z�B���tR�"���S�Y��r�)��_EF\��%�������K_��w�Yh��U�zn�w>���EҰ6� U�x��f|��S����
��$��`�ʿ��j�P�y)}�����t��Ӿ�m[K,3z�I`da�����GwEAO�9F�O�Q��m���01 Wn��� bEԔ���Ծ�u&�W�4+�Wͪ:F��"�oZ#voiB�an��!F��T{�&�n��VLd�����ګ�����"M���O��Fu�?D`��yz���� �=m�:�c��+�Dc�K��L�֑kv�|C�7'���l!l�R=���.��y0�;5�+"߻u�9"?�7_5���A�H��c��^00+����*�UǑ'Caf_񅞄���^q#Icd���n5Z��C�V$Kg&4e��խ2����u�G�������w�>ItA�h��'�,��Du�����Z��b���¸>p?� ���`U���N��7֌�9˙	z{�US�������@�
�%d��K]\��o��Z��pR2HU~���
NG��k��Z3��ű��gRi��5����r���7XvDp5[��k��Z�q��o^*���QJ?���q�Ŗ���6�?�)�I�B�V$������6�R/��-m�/^r[0:K���'�f6�Y�RV�)��9�C�,��= z�I�
�����H��F J��bH��av-�n�H����?��=4��,++���Z��?G�m���l,�G/^������8��n%	T���$A[����{q����������R���Bl���$��S=B�J: lD���RA���V�M���ei�C1H���hQp40mₚ����F_������8H�����	H�%˴h�٧M��5h(I^��6�z5CDP��5�A"���#?'����yv!�M�6K�	KZM��Q��R���Lw ��nN�ӏ��Rs���	�]�i�=VK���Y�'~7K�%NH5���7�1�ys�Q��-IE�Lش)��)_���!H��7������B����R[v-���q�"��M�΋�0:u�J�j���/��Z�S�f�
����P��hjW��<��U~Y���@�f�"���n��UcO�M��7$��/F{�9gB�lb٢E����m���v��3��t`��k�w��G��P�*hw.�&j�:���q����7>�ڑ��D�-�C��+Υ��XԿ���':
�_�ٶ��rj����F%%C�x���x�\����_#a߷Z꜄䏣��E���o�^��mObh�G�vT��j?#7ݥ.��'��EC����������}�n,i��P̑ɬ��(1b�78���fȦN�*:�Y���	��/�$/�����$���skl���c��K$�Ou��uMO"�u�4�	��7t.i7�lu�(Kf�l�6zuL�kJ��H�ۜ$���׃}&Գ:���A�-9˴`K�3�aTӧ�(#����my��>|�����s/�!�b���ܪb�:����k����D���1�C{�Al&*���	��ت@L8��A�%�t��WB���LE�X��Vy���$cQU��"��DV~`���|��zEC��\�����>[!���̍;,��/J����u��9eS�̅k*��뢻F�y{ȥ����c���BJz?w�@��u5���3��~�F��g�obWW��4���ն�6&2���o�0?n��,�`�d�/*�^���0]��K�;%�WM*���p��kNe:O$B�y���/'���a��ƥ����h��KVj	bT��+&C���b}P��V�z��rzf�[�m���=fp��MD�b��f.��SP��?~�á^�i��No5Pd:e<�>_V���(���<kGHʂ٠�1x<@���x!W���:o\��8L�G�*f��Z ��&zO��0��_�,Y2l���2�E&��N��%��!a�dM#��\F)w���e�n��^��P6�C��E�~�P6�f:^���M�[L��%m#�o!͔w���;Yz��E�����.s�M���s���g��H~=��BYdL��ڣu�[t&v�*�U�J�Q6���|�I�a_buT��|چ�^F|�	������|�9��D|s��BN$����q�C����L���z�l��"�)w�BQ�����dRXi�%z�k�+��+1�ڧ�T����,����:̚�H�]W���s@�w�s����FZ�ABg;����bP��K���^�������r_�J��Hh|���w���ݑj�u��^�wym=6�3I�U���	�
�:C��c���{��!/)����/
�/F_�8���ĕ�µ^�h�z�5�M�.��5�X\ j�i���c��ߌ� ~1^���x'�5j���n%���?�Z~���g	�h�`
�`��d%�9��ؕ����G@�:������`��WИZl���McT�?v�]s��F�A~%��W��lJ�>��i�ٞ�r�^!R­@�ևO3��.XG�"����=l�CrR_5�~�Ԙ���̄l�nġ��Hpg�pe��Aտ��rW�#�f�r���v�����U�ǃ�jr����6���]��b�C@Zy�@,���Pd&�p�ZItez�=ļX�K��8ཫX�'#�C��;�EA]�8�uMF���l��P�{�	x�PF���[^ ��>�������>EA��G�~�]�#0�����[
��o����)bPW�s�%_s@G/7 �0��ʭ-9��/�����P�b��|�4��Z�(^��]̟֮֕�ReR�0|�%c�*;��O|O¥<�囎;�o�v�~�5�v����}�$/,�e�݂7͉ʔ��K��jO�z�r$�eX�`:����\q�!���斖43\L8�w�.� k�d�-8�<iV0�C�V�`U�h21��|Q]�숤������(�2H�jfHH^�QUE���7�7@O�W��F���u#����Ƿp������_2)@ai|�攢n��'�U[��՞�j�P����3I�;�0��3A׺��G��B�-��� �Oq�&�4aPd�~)0�ka��-%9��U��#��u�~���(����Р���wMF�9�&NZ���i���Zvc^��K����ʆ�!#b9�:t����1RԮO&�O�*\��2D�O�s�@(d
̲��A��4�m��0�8=z���3��(�,}�J�˧#�N]��}ߟ��h>iG[�� W���o�G.�I���"[��#4q���!�ơA�������݁��Y�鐖X����X��wk{����'~��m��䙺��5F`	C��02I�R�IM	~!bx�w=z����`	�K
+g<r4Z+��O�^# A�z��ot�*є��e^L�|%�|�*U/%�����<��aj�Eh��,s��>�D9��ɨb��)��3�Lz�����,YRZ/7ĭ�����e�&�,?>��XVG��;���_j�!��?J5r�\�COՈG�yW�3*.=p�=�'	n6^��
erNhŨ��4�3�z&�ڶۻ��xf�c-|�S�'��
Ѥ2��&v��Mz���7��] ����8a�VK%�qu`��f��X6>�9/�r��8&�%?�����#vf��ˏ1vj�Id��m��U���j���4�hM�wjD�9(꫱�"ms�$!T���Zm◄�x:Oa:>�LI�
;�����>�i�����Y�WB��רn�ѕ��@yȬ>�W��u��S�o��c*m�%TH�!��R{��馑�-����xJ�:�9L�kG�#x�a�X�Rj��4|��#ű/b�w���K�n����"�M-�ʊ��'��_ץ��?��&�"�Ζ��B�V]urO�l�W~_w��@��nVݷ�y�fh�x�9��SS�oDK1D��N.A�NbC��Z]�vC3���+�5�@�y�)x����<~�RUL���:����x�O�^|E^�-a0�G��}8�DN���|al���^e�Ņ]����E�H���W�Ѭ��e�A�
�ǒ)h�����B���+��c�ܦ}ݻ ��wO�Z�e��3����&~-iEG{����"=W.���7� �3`���Fz��Ke�^Bs�]&�'��=T���@j���A�1�ܶ���[��wE
Ê��a�Gf������-Z�dھ�=5J�J�Ks��7ă�I0ee��旣����Mx��g�oU��2��1a�u��瑃�XH[����{��"�Hvo�>���T�=G!M���U!gqM�2�����(JKl4mQ��P���#Xd�[!�Op�8�V�����[�;�ע�7{��N�h����}?;�b���C*�8�<#���d\MAmh����x�j2,|�`��������Q~(���� �����EX������js:���M6$��,��t����f�.Y��FA�r�^&{*+�:D�z�7<Y��ceXY��&��b;�e�G�c͌�����٧5���/M��Xv�[끗�P�O���0���i��/�P��"��Sy=�Ⱥ<z>_'_�41G���z�]5k�Y��g���+j�и;)��=��B;� <u�wb�(`�	�b���(�S�MBid<8!|���X����=�Xy�(��xX���[������(�d TbL�I�}%��4�`
���?J�ќ�lR<�{8�S�nZ:79��4�c���1.+�|#�s����ﱢ�K�^�Fs���n`�ǨӚ	�8�p��ڋ}f�,�,�iI�k�ӎ�A�}jH�l"~KFi�Y�U���l�E��<�m�?� �,a�gwJC0���A��l>�ow�^�}�n$���D|�&�
�e�[͠}E�����'���˟.=���DT58�IK�����A��w���������3dO�~!�>j��?|M�]��kx�z�缚��- Pm��J`bL|�E��B���3ulI�Y��� �zxl�N�P��҉{ݯk�p΋�a[w?,�!�w�� �U�:�)eJ����N� ��]ڲ��ct2]�
Ri��N�&t�Ķ��ȹo��d�r"h��k%6ż��
"�����M�����+�3��'j�)(�s��s�̱��#�撙,��h�*_$�Ηn�أ�)�T�i֞�#Z�W,-@A
���3�D�4-�������I�ڑ�7��'i�¶>��Uf�F0�|n��D�������_�@�����UМ�Ň&~fN���*��<�k���|z��2�g*x֞ ��wM�,Ƌ�rv��r��Z@��z]���I VTE�D���;�.�_Ջ�в�k͐Ngc��~uC�]�vp��+7ճ
����O��I&��a�?�}D!���5&���֎�.j�n��B�s�� �H����p^�G��F���@��p�h�r����xM9 Y����%Bl�@{Hl�w��8��z���A�4��R������̨����N5Zk#|M���F=
��z�ŝ~<b��<Q���U1�2��V.�S�r^I�q�n� �v�qٷd:y�)�N�GIHO'x�/sNm��fx������ϐ�"�S�m�V���g�MԜWm�F�i����>p��ፘ���#ά\s&����G�Y����	����~r[��I+T��?u݌����l���������V�XE�h�;F[G�p6@U��'_�A�%�&]�u��� ��Q��ʣ��2�*��@o���Hv�[�����r?�~�1�g�+��Z�M�An@YS�u�[��� �HTY\=Ds��\~Y�7���/R����A��x6���#�B1�L�� w���v�)X��'�$�E���͔\f���`��}�>�D�:�ލ*�t4����w1�4��W������3H}�>bR��U�	N���7
Q���,��m%S�~��č��U��)fv�&�Wp�f�0[�;]e�V �;�Oj��Y�,P��ɲ#a�kU�0���.��J8"��?r��R ١�������"go�YH��c
g�'���L�+��3��-|�3�Ж�IU���;/�)o�e�<Rn|N8��-yN@����ҲH{��St�;�oI�ǯIX�5���}�Ee��Iw�<�y#"4��N�K���4�Ҏ�teZ-@Q��fc;e.�
��|�JQw�_���eQ�b�M'6qb{V���q���?!i��22���[���q��63R��̌�+�{�Ii�Ms���`q8^����xJ�S�����	����4�S�b�pj�E�Y���O Բ=x�m�%�;�ir�@`�u��H2�F��� �����l�0�^+gr/gVUgǨ-\z�f�3>�������+�V��j9o&�`S�:��2�#�%��7����2_ב6���M>v�ʃ�V#�R��� '��?W�T����U�Z��r3�K�;�����f��CJ��]����i�*ԝ^�x�z��C�- {�y���~m) _6���X$ŲJ�1� �OB����J���;�s�
��[7�[�ʝ�X2;�OIl�iJ[k(}*�.��u��@pM�3��e��2��"b_�@)N��?x��uΎC^���k?���{��J�c����	nq�,md�ￋa~l?��0 2¯�@�yL������.�7�X���qz��y����F�D���'8�����4b�q����_}ڭ9sM�6��ި?��i.�9NbtX>�lՏ������~�9TY�����X���o�?Vr(�ه�e�{��-b���$�{���F�"(N۳�S�¯Tğp�f��tK�hr��2'���1�,e0<Ȋ�$��[o������[��x�}O%2��:�c�U;ј�^����<+�!�ԃ�G�N5t��~�m8`M������U8ad i��m#5s>�����Q���-�f�Ct���8�'��+Z�j��q#`�y��I0�/��v��f�S���s�dl���[	�c����4N�oQ�?��te5��|�
�9h�좿 72%��5jѩB�l]nřx�|4��p�< )x{����0�*	Z;i����;��D�^[&w����g2���g�y��u���HSb>�mԦ^��=mY��7�E)J1��G�	�7*S/<��}��E�qN�����ؕ�r�&�1N���Y`����j%�t���'If�gGҐ�b6D�Z¬-�:wxD������5'x�"�|��S1�/�ˑťX�I�+:VN�{0�����Q��U/�$�+P���"����������h�+\��*�����X�F��AcR'�Nf��$=��`P{�
F�����Tw=�v2��ʃ�-O���I���=�]�(�t\z���C�w���`��J��Rp� �gx�ti'�؂m%�PD��~cD��n��p����H�v-6]M�e�'.�7���t���x�q�̊1����VzU��goK��ES�.k��=���+	�fM�����;Ŀ��L����8�J�HGH�a����������;�>�Y�i����>�B�� �6tͨ��0���t�g���&/!�9���mbU�3��`|�?��8��+R������4b�~b�!�d�XwVh�Y�ɝ�8�L��}�Nb�ĝ�h�C��;՘�-��_�/�`����&|�Y�'~��A=d	Gt� ��/y(�<��L�H)�2\����MQ$�I��n��#p����|�~�`�[.Ǘꞕ�Ė��:��|���
�IN��lL����\{,];=>[c8�D�l;=�E~�W#�aŇ4�|�'� �j��pR/�3ʿ\HS �����W� �'u��0�Dz�K��=ߛl��D��������"���u�\z�A�]{t�>�4��S3�����R.�/?�|�ң][���XYu�k�@/�l	#�KQ��!���.�d�xy��Q��4����^&(=�5D%��GzPJ�0]&$f�MV����)�c6���v�A&�q��CN +|�,A^�"-�0��˰5I��bn$�e;�2�/�axn�֡��bT8��_����	��MMQ��n�E�9����0��<{:ܸM$�ۈS��-]C	 aߌ M0<-����ޖd(lX�99���gٚ��� 9�g��g�M�A=5�+Zs�v��R|wv�NÝ�Q����E�»��$�|}px�[e#Bv���;�c2�[�r�����Ȕj$�5�y�6=b��p%��/��c%N�P�?P�
H!kxj���9��`��Z�E�>ʈ�W�V~xɃ�D1~S�fY��1�����)(\�0�o̐��e�t��j��G �&K���ٴ�?���	b.��?w�"$���e�%��
"^ bֱ)�����T�U	�m uO�!a�1����!l�\nL5������f�E�4HiҔ3vm�S�r��"-�oL��}=n�
mY��<�GX���,�n�r7G����צT��cM���N�Dx�MkV�i屴�N��,j����O������(a�_l����9J��h�kH�tb�<䱨�[�\��#�g����-����� �4c�)�C��5�f���&P���^P���B���)_���m#_�P�Ŧ����iP���0�3-�����99s�.�{,m�?�o�N�:.��S����|�ߕ��#��4�hc{�"H<�	Y�����$���{Y��º��.�K�&��Ql^(*�'H�j���yI��!M�L��u5��d�#nP��;�+'�� p��.p�Q�Ÿ���\k�0W1Υ{
H�J�� >3�X,�ᷦ��LQ�&~��}Z4��n�w����T��c#jT#r�蕗W��x]�^k$P��B�B:_*�mλV%���x�Tڮx�����2D=�j<�1�-�iC�Kt����H=:��Cb��m���u/W#��h�ݛ��ʈ(D>�i�N �Z0�l|�o���p��T�2�mg�0٤��5�%�|YZ�h��+l�F�Z���.�QDS��3q�/�ULI}�m��������4(�����֌Ӂ�z�7�<hY%	�s'�CA�Y��Bםe��+�gs)$̓�4�A�ԏ�E�R���)���
ӗd�!�ɼq/�J�C���Ul�����R��rD8"0�5��E��Qz�<1M�?dօ
0��8��@ ��Z+=��%�{�FE��~YvJ�f@m_/�x�G�;B�.c!�{Xa��k<�C��N�!��<;��$���w���"9uǡ���0��3e���i����ea�T��A�149��V�
7�]/VHIJ�l�����.{��Lٕ�s�dV.��߆6�Z=W�� �5A��B��[xf?�L����L��v4�!����@]��%@ָz,/
��/  ۷bꧽ+�m{D��:���\��-&�$���[���6������������3:Ź�iukqZ&ݔ��D�T��^�`�n��9*P�<�u��x܎��9�79$>(�לC��G̎���o��+���g1�I=�R���q�<��آU��V�wDi;~���'�ǩ�h4�*�> ��c>%$;��]�q��3p����.���\06D橧��@hH�U��QJ6eN��f�2;Al�͓�Ƥ�p�-�}Д�)U��U!����\tØ��}sz�.����2�ȴ�l H��8~�u�V��S���QA.��-Rӊ"�d7�_U���5;.�����*�"����م1��@p�����Ҟl~�+�cLL!��:ڐ���;�"��p(Id��0������r�DGx���δ�[ �.��]��W���d�Yjd0��j|j�Y(T�X�l�,�v%�8��X2��Ga-��5t	0U��J��W�{g��>��Kk��!�1�r�r��N̴�����i����}����*lM���$:�����7�V�	��4��"Xl�^����$v�Tzo~"@���}��E�ɗ,�LS~��c��:5ْL$��AH�(Ջ�P�њ�[o��.���Kcc��zF��p}�R�ZnՂ�DF`i�OM��3��@3 �N٤��!q��,IW'?F͸�4Ƿ9����E/�{���t��D�S�$��4.�G��%�`��LRR`��O`Kl©1���A���l�"X����$`���z��7�3Ի�q�;`ސf�~�EuvK�#��W��^	L?������x�ʑ�����$dox��%Yr�Pq��V4"���'�<Y��n�=�$���d�g���Xņ��{��Y����}�����N��mR m5ZU��K���Sׄ�y�NHb�s�Y�ԬN���4����Њ�f�V��� N�KzV�VG���)�3��[���D�t�a<�I~�AL�)q��׍<�-0p��)^��k��H�lx;4�' �A�0��eP���.�t�[�=�;[����x�Y5�@�/��,ɔb[>�2�W(�a5u��Ŏ���OX�/%1����w�ҿ�IH�}˶{O�1�2* �u��t�-}�)�#R^��r,�A���e죈v*�:��뮏՗:���:�����'��Z�=�f�-�Ǔy@����u����X��(�
�ADM�����+���1(�	׭z~@����������q�~��a��Z?D!9��G(�!"$���j��T�}x�ׄM6�#y�q�k�N���d�UxE����0���@2�m���%q4��Ppm�E�0�nA
`����� �l,���>��g�9ֲ�K��^��7�/+�_��|N,�?f�_ٞ����|�6 ���9�yfa,t����ɭ>A-6;��9���>�w���t��R�WT��'���P�e���V�Ml&w�9>��5�p~M�=��%t�(#�C̣B,�RG���\�3�`'�_��`�~�D��Ś��dFI|�����������񋂧P�H��Y_?K�x�g��*B�Z�ed��T��C$�)��wq9�>�Ko-l��;�7k����i1��Hq������h|�^�
<%8����W�^xIM?�Ӆ�C���9��Jx���i�5o��0�R�����O��ؿO��t�j���,���K���N@��1�ܐd��||ζz{Ww�l&=L���6x�2ӵ�DMMǗ���,�U��dw��6� ��G9�%I�+_���ϸ�\cӠ�~Uy�~&�V�k�^� ʃ͔2��H�v�$:��tD��v6�-��Kx��kF��r�X��<q"��RƼ�K�c�n�:g����#���#>��G�
��e�2T�s�lJ�5������ϙ�͋r�?\��wl��3;�}��p�W���r!�����[���q�X}T(��4���r�N��2�����<ڴ��b�B�k�]sR�\�9���[�	���ϡ�+s����8?�l��ߴ���޲�~��W�w�ʑ�z�6�� �.�Z0഼�]~No���Qs!1�1#K��H�|�_	d�ҭ���0��4J0r�D2 M�A�/�/��,R����M�L�j5ڹ[��Ϸ�( F���3�Jl�P]�8����`:��������~E���%YG̒F�-��JT��P'����WA�j 3�ß�)�HƒA@�0�
��X��`L �h@ř)�4�d���T*�_U�~k�u��ٱ�4� �8项��*2�Z�#���\�?YkH]m��p��	B�0��뚬g��+-F��/��1��i޹P�[�3�$o�+`���Oq��r3}g��ۑ��ńu�V�?�	"�ͫ���&D�������vA�xc��ҏ�3YҰ�E��U�o�߈�~sZ�Їʝ���C�0n�zN��>jD�}�tI���2��tq��ٌ�b�V<L�`��	�gpM'�|�~���9��)��v�H��!;��O��j��
����i��)�O�"���I��a�`���iGO���mh��g�	��  ��Lɜf��G
��6�p��ӭ#@`fn{K���b���̿4Od���*l^���H����(��{�hX6@�U0�?�q+���%��Vr�1	�#��7:�0�T�x�`�;��pP�XO���p�gK��㮱dѢp�O+ �s/ga�ͯ	,�|룺�k.J�7�h������s�+I�#'A����=yX��,���������b��B lL�$��G�C�%8Hm�?��{}5+|%*$4Z�7l��k�@���x���ˢy�T���4�Ѵ�C�R]k03�YbNSa�韸������8���������̟�=���3��9L����JV����xQ)���.\l����"�
�4��� H���$�	'ԕ��GV��W���1� nVE��A�����`d��S
�:ˮ-K#tz��E���h)���=�:�y�3B8Y���%��Q�&�����"��2���YA-XR�K%�P�ƺ�6��h�}���'eI�o�O�wX�EG���!Q�����:�����z�]�xgV��I�o?)��R�ma�1W��ձDTimG#[�<Cg [��s.��|H�
�O9t�-*g�-�涧"�!.,)4	���Hح����,����/n�Q¨����3�O.�ˡ��G�y�lbp�'�7�H����R	/��ΈￎÊn�ևl�e}g�.��uH�߳u� ��q��$���=�oNZ�+ >��v���%k��4#/�uZ=:�^ﳭN�V�<˒�)"����c�g�q�A����f՟P�6��ww%�Oi�:s���CO}~`tN�k�q��F���Qn�2⹞; �1ou��<;����R������ˏK�@�HXUnFJ�ڵa�.h���%�H���ևD��Fn�A�������~?T�/Y�)�|���Ț����=Y��db;� }�e�])�X[�$t�~>oE�m9�y��L��:0��@	���{���
K<ܢ,��@lnh�bRl-,"�yo��	�F�����K`/�6	2�yL� �W��2�ߎX0��CǼόz��ǎ)��!ɨVC9�]��BxK��^H���D��|D����ǲ�p~��F�N���]�нl�?�F6Z4po���'H����k��P�.���s�+]�Fx�0�pФ5�-��#�|u��塼Z��`v�\��N3�^~��
�.V�����j���� ��Q���J�?��:��N�7����=e����ҟU,�r�����]�;-�0��W��z��E��6$ME���9��^DĉV�S��^����C{����o���1�f�2{�\��Wc�E��Z6�W�DmYrV�p�d��n�����&��Z��ю��D�uaH�oU��b�@H�o�0�Ϻ�߀-��̸��K�v�cP��N�كDj~xJ.�vD��Ԫ���G����������1���t�@��+�\M�g	�H����<�zi�,k'f��=�{�	�8v�ꪚ�w���qJ����2:)!8��w{y���ղ��- x�%�~p�v�H�WK�u�D��]�`a��s�o��% s!�Z�I}=��rv2�	~��e���x�N*�^�����R���3"�O��H�QU�G��%W���n�Nb� ���&5�]>v���G��ِd��r3��n���^��b�J��0%ҹO[����sT�ss�mx���|#�l����	��"{�X&�7��^�Z�7J*r29 �Ac�`��2�8Gw�E{,�����ڽ�/�����7(r�0�Z�&�
���V���H�=����R�勄�$�<]:�"��EĦ�v���Y�ӳ�� K��!W��jW�r��c,B��v8^���􌸡����׵^�U�l�Y�oU�_ΪT���*��p-��Ҋ	^��@��G�e��5FǍ��4J"v�3��{E�adl^Ew��N��6��.	�4�~�X�q��:O�Nâ�>阭�Yh���,j�t(a��<�FN��Ϯ($\ �s�ѺJ0/��d��N�׭'u��w	+����9雊�N�5�.vç[-�.��SZk���!��S��8Ǌ7v����l�̐�Nqa=�-�r�Kn5Yh̻�Nwɬr��<���Ok_@X�����1XQK
>\!�&����&�����Zo�/$j9<��>� ĝ�c$�Ѳ�g$`W���Y��w�zHH��?>�+�c�h��i!>�V��?R'� �B�����:���yU<�fY/<&(�&a�%�����Ä{�O3�
S�!]B�AB���7�{2B<�X�JÃ��)���o@m�G(o��c���S� daWC�To}_������<�HQ��MUrr̆��T����S ��PǛ�J+�����[./{#���F6�H�|�~��:�"1+�=�0���C`"Y�.a���)>)^nD��,��)�1��F�1�!Z�oP������c�d�ke��O�&8xˉs�}�H�`�LAB �Y�M˞o ���liJ�źP�gK�!�Y�d���oR�|��u���"P�����`3s��Ra`�)��,�@�$_��߁b^G,�t��g�x�2�+�BI؇���,2D���(�01>'୘"��e�c�lnG`���Sw�I���>�b5�·�i;��ڥ���催�j��L>��G\la�����뉅h�C��������ti�^ېl�5����X�������w�D*$�}�/NqIw��3Y��Oo�w	�0K+�"�G^�]���d#i}y�G.wO��Mr�cS%�?X���"ʋ�`�l��H�����w��x�T4j��N��H|y�?�>WAM��gN��4*��)x�j�q,�łj�z��m��;%��I�M"8����f%�q+��O_@��6�B�vQ��7�tx�Z	"N�ZX:�=��ʯ-Զ s 1��6Ն+xU3�"�Xu1I��q�ʑ	��U{�)����%	�1!��[��F{u���-���m]�yf/�oZS�D���1�,��m�/+�wOÎf��V6���Q�,`� �`�#D�4j���-7�?��!{3�	�&C�x<�@���4q'[_I����gN�D�w�ǘy"�@M��J^�0s�I ?���r6�Zms�v�;�Ű��]��и��WO�ZyGR�9s�]y ���J���	�}�Ͽ9���_r��L_3�P[��{�����
:&�K.�5����0�tq�����]��{/3��w*yE��e�C?j�3d��K^g�wi�`;O�fb3�S�l2��`ܴۓ\�}0g��q��9����6Kd§Y�/��g3�u���M:��nvSr�Er����閈�zIB�Xl����$��d3���s#v{���t� C�Z����=���ݥ����F8�]���}5�����I?�
�n����jF>�$����������Ӱ�>Q��1��˱8w�SK
D<��sΌc{"p�� SW�a�.�]�⺺�to{;pn�~�(-�)
���v[��
ކ�Iぃۛ:��8�07���_���s��ح%E�%��GW{��u_��mq��MUr���8}�c�I4�_�����Pr���F��!��w�=�(:��m�i�_J0����J�3;�J��� �<�sp>�Z^9�p�.���+��S$.�b Ϧ��Y/P1�ɵ~��DyM�F��N��o޵���[(۴6ͦ�ӽ��8q��~��,�&�;�K��6:р�9�<���ڂ�*�
#k�%y����*�����j���T�b�c-ڤ����&C_��^g<�N��~@���B��|���x\M��E�`��W�8�4�Wh���?�,һ�����}���~(xb�8D�"��лx�4;͝-�'�����g&1aJ���S'E"�'����&�9[/�X@%��a[{�w��(�ڏ@<K:�N���U�����/��d/�[��u^7��;s���/����kU&��8�-�8�����?��L��K	������T���~�fF���g��[��PtK�{��I.2rbm�U>qB<�Ʒ�|�Y�5�C��,��G�Ʈ�o���	�u��~y�����t�9w��q��9�z3������U�����y��w�C�q~�y�ނG%�-.۪���<A�J����Jg��
�h �|�X�n!X�/;�g��'Y�I�S�|�ᕑ94so�qru�g�$CJ���oy�H������(���"8�� m%��W��d�����ߕR�-�_o�
� �;��~%Mȑ.r�~d�g�Am�����C���z*�_�h,�;��fa�[߂
�zU���ڐ넉����o�E���tC��D��I���*'�o�8�Q��R����Bx�y_;=
�Z��1'��U�ź�&H'���S��&L���9�c�����?d-���.��!�H���,/LlQ�ߎ�;��@��-�?r�s�v+s�C��c�up� o�����]Zİ�
�0 r�)vt{h�&(���eRsO[�V!��0��Ū�Xv�Eo�������i"p�[��f�>L��G�Q�������>֋�O�f�7�U��������[t
`�d���k��Ғv^~�T��B�������##��������eX!�W�i\�#��ĺ�Z
�4�U=��[��$]rX�T�P��|#5�:��#"��dx?� �W��*�D
U�t�f��Ѱ)L��fb��Duu!��-�_�bv�� C��Yo�.�W=xwgb���{�B������(Q f��`P�5���3��}K�ư>b'c+bkJ���v�aF���s< /g�P������)c�E�P8e-DV$�-�W�k;XG1HS�֮F.j��<�� ^`���#��'�4i/��k�>�+}kΥ�~���i���8�"]����t��l`���KLd���n�CY�J;��$=g� 
��/  �����Z��!=�.��$n����Jc��R���|4Fo�a���m��<\�\"�e�jj`�)�2��8T&����pM�5�L��-F�Y��D0���ݬD����\��$��z4AE7)�n)�,%���*�'s6s{��q�t��I�}���t�LC�:-��(��h4�*�> ��c>%$;��]�q��3p����.���\06D橧��@hH�U��QJ6eN��f�2;Al�͓�Ƥ�p�-�}Д�)U��U!����\tØ��}sz�.����2�ȴ�l H��8~�u�V��S���QA.��-Rӊ"�d7�_U���5A���vX�m�����ߗ1�49��$�s�S^<+���#ey�j\�-�c�N����lK�T:�{��6��n�I�:Vj�˻A9�|6$V����ڮ����h��BQT��zK�.RE"-L���{�PL	ʦ���hc�]��v|�g�Iv��;���U�>\b	��>��
&��:b�WP��z*����l�q�m�CUq�Ҟ�<_@����@��>�|�|A��Ǉ+��54����:^�<qE'ٺ�64���~)#��2ӜxW�;��b�]��ݶO�ݎ"=8�ؾ3T�jB��咓x��Z4o+"����Z�g)1��nC�ٕӴ- jtj���A�*���^���`{ܑi�@����/���i)�5TL��!m�� .H�6�ig���S�}����^
�9���J�?vĽ�Z�I�|e�w��-&��;�p��;b�����{�H���� ���Y��a0�2�s�޺�ab���M*&5D2C�@�Bvh&6�kH�5�;s�`N��ƾjc|���V�z���xc������Yk�}��Ԟ`;�B���])���ǣ���N�l��sA5/$^e�;\�	J�x��E#���Cd��3�\��I�ѻ�K�TŤ�ʃ���\��
�Y�HUG�Kа���2Jei��T��~<�$�����v�8+~�PG����֭e�yZ,����M���<��=��,ٻ c���U-
��?|7bi�P>��`wb�P=��=�3���g>�}�(Q���~�DX��m�/FFMxا_�S���s�F�; ���5p��4jؐ�.��B�-FG�\��"?��3��O����J��u�*$s����NduXw����������9SID<���#���`�M�x��(r���%瀔��V�5�7��6v{�N��( �+�����a�䠞#ƕ*Hs��P0�s}��ة�!f'pä�[[Y�����:ђu�@IW�5F�� ?��� N���&�I���[��?7����[䇜&��z�H8��֨�e�I�)P��懑��}a�^'�!pz���g+Apa���,F-�#���[�n�t�����f����.O���z�6�\tw�3�%���k �f�}F����0z#�ڣ}�-�Bap!��^ Q�NX�j�Լ��j2Zس����5���Xj�t����W
C�һ;�B�s@�C/=b��!sލ��%�eZR,Y8�N��uw�(���\>Fq����)K�3Nζ�U�ú�B��H���e��4���E���W������b����"��&a4W�������ߏ��c_X7ٲ�PF�v�������?���f��v�����l#�!��<��ʕ��������}��[gf�팴�d����?K��"���lG�\Rj]��.|��H��� u��J�f��Thu� v�d���J����+#iC� �����h��K14���	F�}�����_�\(��(�RGl`%�jO�!<���J��W졑M���ﯷ�M�����eZ'I���P�\��2���>�.�]��Q���@WĹ��{K���u�q�j� ]."Ƴ'�r�#R���rv�7��dfS����E=����6߰��+Q"4�=L��{y�oQsȭ��T)ٕ�����;ײ�X�-@�ξ�F��3��h"n��-iĊ� 藺���9����p,����Ţp��2HN����^}�ѵҖrC���A��o'�`�!�����q7�
=q�U��h,_��k=�Q$�J�Å���n�"�<�b�|�(ošĿ"P�x`��~�uG��.ջ�{b#M�s�v 	�`#}f�I_��H��4��W#u�1`��!إ��6�D8��>u��G�!���tA���aD�i�2Ģ�e;���q�bF[g���kz�(�/���Hj��0@�#�P_�/I���CR��>đ�ʎ٣#Q��mJzmŭu�K�K,cTN	d�0d<wf*D�b���?��RMF��rF�mdk����U|P�>q��8��B�N?Ѱx<��gzΆ;����p���.Ç`�����VL��1w1P�����j+���!�S��>�8�.w�Օ�rSap�����k�yE��ң ߣ�T��'k=�5V]��id�G��^�E��A���H���U�q�Ge����&�����Rn�>a�R�ݗ��2�O���/}i$(u�a�L��^B.��Û>/�A�/�� ����"�֕�B����7޷,��wXI?�1���Эo�R�UDnP���+Q��"�v���_y��ҏp`�)���:	6\gp�� ��/�t6��B$��Z�;Tg�E��ķJz�`aH�e`3��
���̖��L�_V���hfp�>�����bS4o��/0�� �H��^�!�S���C(d�f��d����EO�4�i4��}���3!}����r� KWcz\I\K78��n�n���պ�����'T#�8�9�}���r����.���}����#�<ͯ��m*j�XtG��>�5l
D��L�H�-H�#zЩ{پ��z���ѕ8������޲��p(�\�|��_n �#{��B����P�HPB�6�������2ܳc}����DUH�w�x~F�5�^��IS�����,�%�D��m��>�j�����
�W�l�3S/�,���#�nX<���g����Q��L���6iq��3��X>�a���a
���R���Z���=$V�Vi�k&����)�f-됋���.�H�f-E#��ASS�_{vS�;��QDY_y�Q	�ǔQp�飐�^���$/'	RjޮI�Zl��*2ϥfS�����y$�`��I��:Mϊ���Bo�"LA'5Ay�������
pVbFID V>���eZ��]�Uzgh���FJ�������6t y�'��S���WV])W���&�?��Z��s	@\0�"�.7��F���:7]muyp�O#�p *~Er��k~"X���}�1ǔ�KNm�pusQ�&Y��|,�[6h�5�g�lҺ�	͙��c՗���"nrz @�Dp�ڒ�
%1p���Z��Еwv>ɒ���^` �~0r��,��̯"�ˉ��n���r<r���/�g��q\�?�9��J�)[4D~�Y�Q�}p�LE�Z�0=��N���p��*�S��b˩����e�<;`,M�g�sg�xw�Y��A� $%����Cw?�:P��6*���ҏD�(��ͼ��hGB�v��gsb��/�]{(<o�;�x`�vt����ii9�5紊SX���W��Ϊ�^��Q����� ����� �я�ܞ��Sħ���1����D��͹y��_7a�T��q�%�{����G�(�ʸ�=�^�Dͪ�5����QN��:F�\*�.�5��Z^��7�阌 v�'���J��&g���R�p��!���P)���&��"l��G�g��Tn�`Brm�S21����hݖ�4��'���c��ht;f����t�rC���[���}��DY�S�x���L�1�V�,�����k�Jj�`{fx��s2�A��x�	�B�X�j.��:���=�m����p��Y�������:�-�M#���9��Y멷��#�����B�a�'ᐦ|��J����͊J!Y�ӸS�3���	5��C�F{��(��-�M���`�&-�W�M��fU���|U7��E풃�J��'��8��u('�W�<��nG���B�n��+���0�ؚ��&8�	�fj<XF%�J
k����!����D��ݬfN���v������قw���-~K�M
�@��C��(j-M��X��E6�tmS�p�3�bY�I��a;�c�&]�g��ۅ�q���h!�oG����f��@v*��[�U&Su��V�B9�>�J���� ��@π/$C+�[�N��Dac�#��)^���1lV�)�=h&�����Lٕ��s��Q�͌d�D�sx��3E�nFpq�.�D�11������/��x)W���T[��P�b�e�`w�-�jrm;?zn8�g���v\�6ɀn�����^�49�NQ�#A��B�������x���31<�ܐ4���6��*0o�|��Ȳ"����K<G�B����V���W���1�8d}�a\~��K=>9	`],_6�3�_O�\�� ��X��<�UjE ��`�`+[&Y���-b���.s����3��8�j�	���J�>l����������a�� ���G�x`�¶�q�}��0�͍�	Y���9�[Ɍ���b�	y7Q"OCw�?�9�"�2ՌD�WRі��$7DŒd���&�華��W\����'�]���o��*v��T�j�u
�J�7�"�F�����
��>67��8v�^p��2�i�o�τR=�pҲH'�a���r=��DR����-l]����[7��֙��C~�S�܀�r�Թ��d��.���8����|FW��`��vں�qã��g<�?V��A�ѯ��~c�ɛ8����y#�?#����Xٜ�.�Ԭ6V����:=H����f�yQ�Z{��%�$<0e�ꆜ��{r�$�Fg󖓜�4��NL|�j4]���4u&��NCGef�+2��/�&'A���E�^��L��4	��8��=n�>B�BV��0Q�(�P嫝�*����W���u��+i��16�O����Z��b�k���Ս[��+�1g)��K���=���2=/��%cı{�쓭\�_�-Ċ;闭b�y&���3�r�J��r�ov!�Yz&-⨲t��O��}�x ^�~��B�B��*��O>��)»'��P�&�`<��(C�p�E��-�4�����QxB���ZS�uK��cKl�W��ܴ͸�ı��[��������=���a��U�]ey7Fi���T��4N��0��Aϰ�������Py7�m��W�½ tj�k�Dm�@$! �I��
A�޵��Ff�8KU���p�N�@h�3y?Y�Ww,�&(�qd��c�K�B	>TL��wo�2�Kna���a`���W|�o>L�E�b�5��� O�\ B��[�͞��=#��_�LƢ��y{�$ �������ҧ	.�V�6��*HA�K|T�e�Z�La�a}{T����-^�l{�6H��h���Z}��|u&��"�p~��1f��ySE��8�Y�v]}�
����hG�/=}/-�x%��<�mu�&~�����t&8�����^�=�ך�j���y;0L;�s�a���p2x�G�b��w�?+��{�LsrU�K&��rR]a��r"
!�	�O;�}�e�`j��4?���a�\k�Z	�W�)_Tj��� ��I��X��L�ᴴ@��T�э��ψ����z��TbW	H\&��e�wh�u��$�T����i�]a�z�v�]/����Џ[u<��e��>��9�vy���F-����cu�9��S-
�7C�E?��T�02��%�C�Lw,��R"!M���R��n�B]
$w�V{+cӰ�)�\�L��CN��S^kzE��œ�T5��".>��~3/��[d^3ԙ/{ѳ�v$�8���xl��������*,@��o�IP��H_�:��sow_�����v�F��e��w��GZ�אt��I�3��������" �Zǂ�K+4T��V��Cd$���R�8�4y��&����֘� ppY��I��v�l���F�0�_��7�\���+E�o����u���CMڧth�$7nK��^�-!���|[�^�*�	^7t�~�6q��u��m@�j�K��KA�|���XM�W1���Ao��3mk���)�O�`�c�\*�9�B��#ߌ$�Hgi�6jD"�T[��j��Ŕ�l^j�.hE�����\����P��'���Qӿ����'�p��ˑ�ƣ����`o���R�V�)��89p�N��򔌒�(#`�+�y��+4&Ç�G��	L�!����`_���D���)���6_i�`)6��Xھ�?��g���i�/g(����A�=�L�u���X��D{�v� Ǔ��
a���H�Q5���g�����k�u�B��߉x<j-��F����w�*hI���!�՚ڗN�������~�̜���ڍx�VĆ821�袔y{�2�[�۸�]��œPE�j� nHȉ�xP�m+{����7��������C��1� ~�T���wb�<�)��W6�G��:e;2�]F��x���C�����;q�g��Ȗ ��r0�?�����+��P���n?L����7���9bn)�\�S�π��ꢠ�� 'qƞRG�d�HQTpi V�T8N�������.-t�� �hvbw���%>r6{�sI��F���A���+ۈJ�K�����<o�'?
[�c�<�\"�5	8��N�ǈ�<t�0��,W0.�*^T�ՙpZ�1��5(�eApȒ�I9���w�Y����@̼2(��H�c^�+%�;�� ��&����9�o�Q�jp�1����"��ű�iL�ՙ�
Z ׻(��X�VT�g^hŢo�,p�m�%��5��_�k��_"Ԛ�*/��[z����*��3u����d�������C���x����蘬d3�C$ZGk@6��(�bK�UTA�H��M^���:�H$��&�z$�k�e_E;���$Hףpb�A��/�X'<��!:}`*�,��(i;rn����g�g)�dC��bj�t�"AB�2QJ�2tL���u erSf
A���6���M@^!j�m���	��9�2��~Ϙ���څߖ�:{O�̞�6���ʥGq)��mC@)��!0v�y6��#�sV�ɒE^��^��J�Ϳz��$4y`�(����]|!��q}+�������w��?�M���qS�Z�~H7�_�Ne-�(���<�KPFT[%ہ_y6Z�oJĻ���8�����	�s_V��� I�Qq�d�l�����[`�=�]ܡZ�Y�D9�/T���t�$�D1D�A��\ ��d��I�u$�v���aC����� ����Z^��.���G�q�m�k6Fk��n������ħ7�H�	Q�Cņ�V�46�g��$�t����D��yl��Z��9 ��GN�9_|;n�ޥ@����#�U��U1F?)>)m��7��*�q����˕V7ͥ"�hF�����+�*���=��=mT0�3����Y�����/���YI�l����zR�M��=����a�a�+�Y�m9�0cЖ�Ө#g�E��uM4n2�U�9�aM��0�r��G�$�z�#ŏ�T�:�W�,�Q�4ى"U�o�B�V���0��gq�W��(55WwA`4�9���zz���5��j.���MSW&*E��b�$��F�w%�@aaC�k�D�M<���ã&Z���n�@}��e��ʐ�X����N�?E��t�M��&��	��sAxO�M�t����%�[\U�>�O]� 7�O�׌K4�r�=���Ȧj��J)��0�g���QB��(?u^	-�9Y�35���HXU��П���GQJCW
�"m+v��4�9��F]��K8�O*Ry����?��D�p�O��$���=�W׵����3��4Trܘ|x���:ְv)�"4ɃQl�`'PYPIt�%������dE�aӇ�v�y)+�$����^��9"u��o_|����]»,�q�N�����
� ���Iz���n�:��c��Ξ��6k�xs�(~���
���.Z�7�݁�r�z�fR%�/^�C
}�(v����u�}� S0�y�=�gu����GK'�iE)���D9�T�w��o�V��7�t��Y�0��μ�n�*�yY×)���Q�L����S�ؗ��������2�$��L��xśvN&������1;��M1n}����>s6�khior�^�����g�q�/�j��x����C�hoHR-��;����>���`/�o̍ ��}F�cϽ;��$g)��
vohM޿�V8-�֙Ã��/	��X(��X�tE�.�U�b*9|�4���@&�l�����8��Y���K�EJG
�L���A���[�������=Kĳ>��f��.�Ex��~V\&E*e�����Z��'q���;���]NT���0�0w0��xD������K��k4E�ޔS����V#�����Q�����X>��+���5���d�+C�^-"$�{M�3�]k������^��F��	��F���l���ȹ����M�K�N�8��bS�Ν$Vdh��Zw"�	�sP���J���i�^|W��K!�`q�Ex��+E���=��V�����̻���)����w7P���M���3HMy�& �
��}Gb�}�%i��`{�XD9�o�u��o����+��>$@Io"�{����0�t#��h��x`���_��m�t�+�F�Dd��_�V�-��LKq��bx�큫�A=�UT"Pg]`Kr>a�n�G]��T��n��߼�y&!��-;l�C��� ����+���h�Mx�X��ciH�7��R��M"�ԛm�*�CÂ��d�N�/�}yɭi:Np�ǥ�}�ڧ/�R� �r��w�L��79�E��L�js⮀)�z3�c%w�wx�����2��^�(P�Rщ�B��2��j���r���V|��=�
�C�ܲ�I�)B�W�P�F*ؘi� I�M_�9k�2#���˹=�*��w�?�����V$��6�s9�OxkWl�i,;�HUzX��B$��d2Ə�Au�Ŵ@���'j�6d�<�=���_����`���y��h�߽����c{ǘ����H�|_�$��풳F@�B\)��c~�˚��E�_��z�y<�&�b@��Mޠ������J�d��i����eL%m��Ϳ'��8�t���]4R�>�׉��:��܆w��$��Y���:��mMu�W�6� 0��/
�&�Z�($�x �|�B�,�#|J���_��85�KwϦ�}QD�iPu�9�k�hU^�K5I�L���Dn�+e�x�!{��Dpv�� �	tCp�n�}ߵ�h	�������&1�ªa3�W�N���ICŢ;oV�K$�UR7�d.M�mִ��|X�
k�BU�����߰���3Ӌ��X]����#K4���Q`Y<\;_9?�mV���??�\�_����oEb�<���V�Ӌ�M
��Hs��md�Ww�%�8X!,f��zL���Q���_�ԣ�>����Y��-�yŭB��R���;��~�t��5I���US��\?�B�tѾ��=��і\�#\�������Y�j�tV#~k��s4�Η�_=���Sa�T.��d*�Ț�-]ٙ	`y¾'�>짯�d!r�7���]]�ˍ�Nl1:_C9�߱Re�d!Ǆ�:�#-4#�:!|;�u������:$���l[����R����0*�C�ݘ�����A_��
�l�ym$�aL�q2��u�c�J�(��lUF� 7i"�,AƩ��&��F*�E*�
��a�@�d��W��ay�x�܍jI���J��UgC�<h�� X:��܆��n}�t����kilf>����b�Ao��/�݃�:���(~���	�W�T�V�%t_(�f���߬&.�Rw�wE��x �%�>X{"͸�%��L
�ʱ���w��J#�Sy�n|{��D�����0W�H��g�9:A]vNK�UM/���*�%o@AAJ��%��(���� +]�]BN�ԅ�t�����I8��������Ye�"ؑ�0|��dS���������%8�YgP��@��X�����~��H�*�K��N`'�w��N��Z�wm�&Ms[�^�=�HT��z^L��%���U4fGddeӻ�Z#n|�uy��@��g"z{j�Q�R����fd�����ܿ�����$�Y�Y󶼮W[�j��-@�jxV�+e���kLZ)M�f��H�Vf��z�g�,!�@��G��6�;�O��CR2���S�u*΋0�Ŭ�"l����l�PV�O���\_찪B��4�U_}yN��dF��o<(.�՛�; +aLU������o�Uk�c�R�1�C�𭅼������ E�4��@�+���_�O_	���ܡ+�"�Z/;�¨o�%��ݼbo�_�V�{j��3�:��%&��_�p.�!�ۙC[<{�&���9�Z�C��y��g������a��i��'r�q�jX�:�y2��[T��O	VW����d#&�0�|��l��u��5R?j�"���z]>��?��NY8/�0�B�r�l���2�k��A���a��W�8ZiW��Y����K Z{����R���q����ͧ����NN�S Ap.�:" �BX�� p��bьo#OĿ�ʦ%R�Ӫ1�hЩ)a(�� Im֡�C�K�ng6)<��iم
5��q�s@~顶U�5���i6Yh_�,�TZ����X�����wSF���3:4u7_i����݃�<�,�؆�C^
���yF���9{gX�a]�������{ʉC�x��+'���ɷ�
���L6q�>;w�
�V��΂C&���U����]fN���M�i�=}Wju�l�ĉ�ᜈ%�*�$��8��\�+�Ȝ�l9�q�[��̘Ǖ�����>よ�,��eE�x�F�pn�?�����P>��v���+�"[�h�d�S}�������J_���P�_k��y���ţ�� IƖ1�ʧ�6T%h%�o��d��X�*S� �h�[Aw�UwI���h���#gr���
��Y�_5�G�*���;���i��%���w=J�b\��EsM	e��i�C�7��6��f�1צ"��Rn��#��,�o��Z1���+�8���v��R��3�R7����uw��t�BۋA�����a�1�l���wE�~9Ȯ��+E�����7�E{g|�+�RZ���q�ꆛ�V��:U���?Ȩ��$2�
���#���d��f+l;N��0y��L�1�ೈW�h�U������c=;�.K��7p`r����1� "��t��p%Z�e�K&x36a9 G�v�YlY��AB�G(�-�?��ȁ�-k};����2Ƴ۔F��q:��Cu��!�c/8Ǚ��u@^�Л�:PC�Ud�Җ:T�t8���7	K`������פ�.����u�OdX�܁��B�%�E2U^�jmR8Î����?
���,�x�'AYecP�d?�����FC�1���*?�vQ�L���q�"�$����پF��� A;��/�	���n��݀,Pc�p�@ƕHo*��S�.��)���{���Ť~I��
�V���	��`3m~��]O'�u�SQ:�4�0D�2���'4u������IXZ�Z�L����R��L8ӑaVqΦ�����M���Jt�N^c��K����|����lÈ|A�Yנ�ۘ^�����x���l��;�^u�
0ߨǰ�C�yt��\_��GMz�"h6���ǩ��e��_���2:�o3�GP'LL4�	�N�/ڒ���K�)G�`+(m���F=M5؅�S�#�nɑ�w�jN�A�j�����;ψ16�����LF׫q��d�O�'�X4�$/pP�39dkO8Xa����>�I�5EѡT�[�E�������ؔ'B_���G]��tҸUmS���V+����5����O�樴ω0�(����;��a-'��=Pu�t��<����w7KP�w<�>MW}0��d���㕃�[� �N>��my��"[�#^T&uz8�+����s%�]�APP�d�d顺u���0�L�2{
���]��w����^�zXf<�S�����(	�u��
���H]��X��2���a�7����?��|�7d�S��Dl�$��pj�^��}�X��w ����y��%����Ղ��˿�����Q�H$I}!����0���Dq� ���e�X��uj�s�o�Ny�Ҡ��l��E��	o�5#�h!���+��������;�;���p?}I�\�M@TK� ���Ǜ9�I�W.�!��_'�6��"�|B:�[�z�ɷ��S{		��N΍t��_b��T�#�W��u������^�8B�sOr��+��YI�l+��O��P��
+��6`�#�3���q�q:Kx�t�B�Wp��ɹ��3"��4�O ��G�л�t�i�����^��0��0$�E����&4��bw���28���n@9���>��u�Y��M8м��j ��L��u�q�2Jԫ�Y `앩B��^�W~~�"Rl0���U��_��'�Y�;�yf������"�l~����v]qcA�ͳH�-��`�@8��0c�9FC�V��s�z�ƈ�V�����^�ԣ�n�y��n��.�Ъ�}�%���̷�Jpn�j��V6�z����;=qI^������o� Z�}�_�D��Q��^��.5����;��ha�rG`&�z�iD�[d�ѿ[�te��-���R����o��}��Q>(b��La���Q,+�O
�Ya�F��9�<*ǀ�����$���W=0����0rfsq=m��N4G�� �����!���)_M{�uҤcN	~��WW�L>�/���#f�Fg3�RZQG�4��˭-WZ���l�RL� N�����=�k?��%��>j/*ݰ�쵊�˰lOC���~�w>>��5��E�e.<��A�-�"�^	*`5�%��V��~m6�L;i�����XK����y��ѻ��U.;Ǐ�PwI��ӝ9\(�N��.$��#x}V�K��B�p�M\RZ���ww{���.�Ut�64�䝟� �����02�2�yY���?�!�_�`�[���K[(6�Ӷ���3f���p'�὇��@a��P:�rF����8��M�h�Kj"j���J��Nƪ��W�df{������VF��xTǂ�W;!���eB�1v3_V�݀�Vpe[�W�H��1~������ȟ�B�U͑eSϝ��ü��.���ݰΧ+��rR�x�T��%7�l֖���a"�����Ĭ���TQp���*fx0�E�=��~�Z|)|,�I��+/1��m3�XIUp�-��}���Bx� r�$�������CS�\B�~~�����![|}�<�u�q[�!_|�^���c0
3`�h����A-����5w��9���Y5��H|�@��]�oب�8]��B��bd��7������j��)�
MJt��,><F �f�,vK�q@�۵� J��셙F��Q����9�O2KUtZH�sS�Kj��2�݉lk���'��:�f�f\Y�K�(d\��J���.�8��-BA�W?O2�f�fjŢWӨ�j?��H6�c]-U����,?�/%j{R�7�G�+���x�ف�v�I���(X[e+�U��z���>���!���x���ZWK3��KY'	x6� lLK��Q��d��@`͝ή�$>Yd��;�z5*�Wڃ���r�1p�>���b�务^�&�_���S<������KnÅT@Xa:��wF����đ���^�,ju�hS��X=���N�hx��#�C�	�C�{F��7+�u=tk��Y�[�\�ÅkI��;���v#xa�3Br�v@ѻk�eG�̀����κ��0��I��=@��Da�#�WJ�RY������y��b֏w6mJG}�5n��rn�+�o���1����3����6{�ENh�c��_8�פ�A�&P�NɴZ�y/`U�ɁD𼷁�%��z�� �s�o���q�<����hX�0+9��<,�_#���^g�q�:�}�r��/x��ߣ�dOc$����AE4�)�
h��K��D�%J��XFe g���o�}����4�y)0��Z���N���O/�$�C�ۗ���8Z�!���o�p^:��P䄇#e��-[b��D2��˂�ٲ&eHf;�ز��bjc�k�?f�w �}���)H�}"����NFj�b�C�h9�d�)/���c�u�t�Ey`�%�[\�����	p�	A��ĵ<b.�X膡���k�4��y��r���s�ULr*h�̞���uy�褞+Ũ8Y�����35<�w�)���;��0��_�\��.�L��]��5����K�n ��>��Zp�a7C�q?%xҎ!�0W��zmF�
��ڧ�n��'�I_
@����\}�������9}�ZC�F�v@����Z��G�𓍼�.�s4��K!� #��a�Q
�Wk��^9��lYgێ�`Y��i�(1(V��9-���2ب�SˡI��1��,L�b�\���M��V� ZZ~m��s�d��{��ұ�Ƨӕ�Eהe�V�}a�E�k0�����7���n+$�F�A�_�\�A,f��O��6�@ı6�ʯfƪ��6�;�J�����Q2��3j�^t�U[�h�����X��Fwa���@1l��v��e4�$;.nc૶��?2[)���Q̽�����]��g�J�T��;����Q
���	Wc+7�or�_iZN�{5��+iQ�Ƒ3�j��$<2tc�r�����>T[LB�1#=��T�ˠW�0˕�3՗�=� ��ؓ}�ň�6�L���ڏ����+�[��ߟC�lӅ��d�m[���]��6z���j�F��g��fD�aV?��1`��+=��Krԏ��lzNK��[~9뉷säCf:��nGݴ�f
d�]Pmww>-j��T˶��8�Lq,<of|R�oǣh	�݁��ė��OC��������tC�E���M܎2�\���6gHD"��0f	�,~��/'���
߿[d%�2�ԣ��h-0	c��n�P &M�+�j8�g�SV<J$�$,�x>�2��E���J�oEJ<�+��4ke�pұ��_���/P��F�I&��P��NzZ�����~�}��p/�L�N�L��(��,�P�t4h7�Ǆ
Z��d��ǧE��m3��� W#Q�� �B7����VC�k|�{�������{7���,OwGϗɴ�=>�O��QM���MK�F^����RsC�7�� r�,�.��Q۵M��qZ:����o�A��j�_�X�q#ʧ�\xc4G$M
������Ա<�-t��W��:%?�2�k��@AWt�&�E�A�m��Kz��g�E^3-��UQ͉�����]V�a��ً9��B���}���J�</Σ������ާz�EbBR�C�E�%�G�4	#�`����.'�8L+� ����g�{[J�r
]�R(�T�A(�5�]V����r�{j+�N�f����:9��?+�B|$8f`Ǣ�!�26=F��:�A%�b��\�ݝ&	E�hKL�}�2�DNB<���;��y��5LA.LS��F	u|��o��^�"IyCM�;�:92oLmد�,$�dg�6�1�I"��Xxq�yz�3��%QDM�����k�-!doD��a�h=�&��;���H� �m��<���<E� �j��V�$�тռ����F�ֳ�pJ��]S��'��4��ӝ�J�W��i�]�*7s�8�3����􉐺�`�|-��ù5N���u��U�s��Ø��,23B�z��땗���x�^R�<�K���GOv�h)���L5UN������*Pr<T�f����P��8�?u��\�֠"�ۖq&ܚR�ț�[���-���^D��2�?JeJq
�]$���S��7��˜�k�#$�8B3�*��&#w���� �� ��Mϖ�H�.�*�[cP�4"~fR����#����&1!�P���r<��i>��=T�X����+ꩲ�1��J*P��@(����ӝ��G��n\X�S��-�>.{���5�ʷh
����'���^;���O�Q}Rf%��결 
;׆�������+�~�F���#�G;��B�7äWv^�}���>��*R'D�T6���t���qZ\���<��hVm]ոS|�I�d�X4��(φN$���<.o�r'P�!\���f=�h=:y3�@s�8ɗ����N��r, ��oy5m�Y�?vԥL��C��f$����A���T�t�������'�0X�����)1�5x���ؠ#XHڪ|�]��o�Ѧ�zu�P9;�f��]��[�%����0����7� �:��T<�_� rp<┞�"nm���(��= �^;N)K.V�m6�"�jO��B�t������0-�A}�^H�����j��mp6��&0��V���HS3k�eWl���qV�������/5d��kT|V�Zi}����%����Y����_�8�m�K�}�-��2�r��e�C�m\����B|�#�GJؔ}!	�hЛ�g��Vn�J�1j���M�_���uK,I����7z�)x�0�0i
i���Љ��0�*/if�n?v�!�l��8�8]���,��X��K����������Su�*�$��?Z�y����nw�w����n�����bH���C��'��f�>}2�*�C}���'}���7�����U'`��S���}����T#f��E�9[��7�w��?��x�Q2�����
�R$�?�v���gh�x��G�OD�A��ְ�<C����Hal���RDh;�y�*�uP�����M�]��\(��{N|��2��u	]����o�߄j��vo:�Ļu������؋�1M%�v�y�G���>�k_�158	�Sv�[�4z%��>����N��Ys�jaD���͎��t���:�t�8���1�xg} �q~,�Ky�a�$��U4C`d����B����3I��	�O ��Q�B���;LN��� �c�LJ��������'����Z2�N%6��+��MW� Wa!112��"b(���Չ4f���H�F��2������'��o�i���.XȦ V�fm��딻�"_���б��n���<�|�a���pC.5٢�� %�{�~�=[�_L3�����"�tU���{1���v�ۖ�3�����3����R|�.&s�"ݡrH��� �f< ���:M�n ���S^�TA´NH|��d�(�;3�Ry�n��� t(&�G~�$�IKJ̣W����u码؋ V�}һ=����d(�O'�����Z��h��� l_�mc�M���V{�m�Y��������I�N���90�/_'��.�����L�.�rzW'#X���[fI�D��>$tb�����<�(Q�$p�{��Z1��$N�a���U}-4Sif��_��Ằ���U"?S?Ґ��YϽ�#Y�X<yv�#����妅iѢ'eM���͏���w�k�Uٵ��7І*�dI^����f��nD�;_���q<,�~6ҟ¡S6_�w Z-�Ԇ�JmbD��X�1�ù`���{U�Ů(qx��=���F=KS���fꪜ���VMl$���!����j�4!#C
i�rnY�~��'=;c�)���Ƕ��Ԙ�^k�GA��RC&���9���UG�}�ߨɶ%����$	(�sȎ��am�%=�{�����6k�]2��n���.moq�!��Qspk���I�rRKHI�eKn~lIg�u}\�_z V������{�K���O��uD�Zioz�K��{hM�����FTu��i�[��-�pYͧ�6�C/Qƛz�����}�]"�dw	����`F^�ȁ��$[P�5�|����ALuۜ�E�0��S��X�;7�A~�G��~��UY���o��ߤD��?a��IV���-�Ԣ�7 ��/A������
�0�T��W,jI�vSΧg�j��.�^5�(���_�U|AX�����N�/_�	e��	�Y�8�7���EJ�WX`��~z�NF+���NB����y��JP�����TiCk�~����.8��B����|S1a;�a�7��� ��i~� �ˡ4�4��
N5Ћc�X�������Jy�!h�}IխN�T��CZ�rNo���c�Z�>TKõrL�H����aW캔�C�[�L=��(N���e��)F�+�z8�h���43������ɫ���Ƶ�� �/�Q��\�!e��v�%O1a�6���:�W+�"ѰE�7���%�uXf����X������[�ˀ\��]��H��Go�.�eYE����l��!AO�� -w�����
��;7m���H�p��2�ٖ/c��8���8�,CC���Fd�Nb/ܶ����!��
�V�R����WؙN�����.�j>�:gڷH���Lk��"y��6�g���9YN��GO�I��Jsa�mWH#���Q2�\�=q�B@:�gǘWW�"%T�_�L]͆�
��s�WEM��m2�L-��fѲ'Z����Mv�G�7MHHӟ@�����_�_�K9Qt���;F"��p���X����>�p�kUԘ�;�Y���J�k㵣P�Z-���B̝PnF�븲<���p3�	b)}���-�9Ճ�&�`�W�<	�Qg�K�C�n�4��)�?9�u�n����&I�K��A�|�͋���m��<�(0%��f1�`r�m}�����aO;�.<)�����R���|��,0GX��Ϯ2~f���ӭ��Vl*�'L턋�Pw�z��&$�Ed2e��?6�Iv%i(�q���I�����l^p�,7~�Y,�x�r7��O/�bv��t' }�2������$Qjs��v�~j��Y�BK���;i�������H`%���jk@9������]�i��O���!h�X�������K����
M���5�SF�Ihb�~����ُ��Ƿ�G6G��5�C���;�af���9�*'cw��]Z�9&�g�_���s�^jTM�t|<���:����ű�|���gDN��������b�:��!�V�0���fu˚�}@5y���\Fr-kq��d/t�l�T����EU�Iwb�u���D&�~ԓ�e��':�/>5g{T�t���<����Pi���9R�T_+���bMa�E%�Jx8�\$Jb� �!�w�ɲ�\�/�3�舆����Sn[���k0�G�Ĭ6[��	�h��{�^;�ꯩ��/ʁHe#�[�!=���g�E{�6�$y6�m������Z�n2����(w������4|�.W��YT�l#�$�w�����"���O��+"���i!�9��.��ɮO���~Y�s
N�<V3��y�mt������D<<՝�#7�z�0�����<�%�����1��>=�$݁��C���s���Ҁ�����Qb~�� ��Cٶ^�I�;���8r���Nk�[YA	0+��\dм&��1��)ׇg�����!�BiZPM��X�jl�w6_شxmX�,�+�SX��Q2��!ذ�?*�d����w��<�zZ��n�=5X.��u�D�RI����F�^z{�|�ל����1�H�Y�Ǽk��M[�;(#�P�x�G���L�}Y$e���a�V��F�=��s'
��Y>|�e��&S��V׬ޔ
���8K��\b��3�xN.��^+!��ܯ�Z CЌK!f .����2���YD�u���9�DbI��$7/���?uq"�S��~;�S�9�SOP�%�ַ4�\�)�5�����r�]\�� K���<�ǩ:q ZnlԼG���/��27M��!�d���vL��`��+�r?���[K�
q���?}�џx�9fO3*��gu� ��̣*�P���]�;�*6�<�V����	�&"��먌\ni��	4q&T>e���.�0o����&����ȸG�����@e��s�	� �����T�+i7sB�4ة?�p���+���~b��_%�y���%m
q�;q����	3�[��~ֱ.����1O��o�μ�CD+%��Ȇ����.��{�lH�QiS�8+A�����n߽{zۍζE���⪒�}�n'�R��5!�.�o��/�`n��t�/\�Z�?a�X�v �m�R0}?��� �����0����8)�����H�м�PN��YM�$&�>K���y݇��i��<��H�Ut(��樜?4z챇PS�+� �a�!S�a�p�P�rX�r�m[�7���F�g+�F̎��e)/�4�5��?m�
3$<����_<o�MW@,^�t�麭� �~mXL]��N�^g-��:U��6{��ڮA>P���p���E8�O�WY'���6X��5�0���!��X�Y.M;;�����HUT���-�Cp6��q�"q8s$�F�e�X��Q�z$`�tUQ^��Ñ���[C���ǁ/Vs[�1�V�APĳ�h��p���"8N��u���U�I����,N��6����J%m��:���zd�ќ�_T�v&$�<����=~�V��|�'�I�k�1t�{�?.4{	ʬkn��+�)����fL@�F���:�`��,�q5�;9h��!1�A��3�&G�ų@�:7�	.CF�p��r5 ,Ty/U��-��4^�t]�#��s����!2�Ȋ.|YR&�_!c���Y�3�[��h�U	y�Aa�,cg�Y�[=a�i�|�����_xA�
,+ b����sXm�$�k�_c�^A�i�58x7���7kW���W��~p��n��Rn>8, �=`Y�ʼ��2���-����wQ��T/��H�&��Z:��;M}��!�������ȝ�;��r�Q���9�#�/�	��9!��Ă�<��p:��b*��2�S1��V�>�:�>!ŭ־�Y�������wh}1��#-9�����~����eR�)9C_����%9�&8��Y�f0�V�m�� ��dA(x
��:'`�I������r�耎����A��w08�t�[��m�I5�T�Rn7'&�� ���߁�_�Ɔ�@�b�SR���V?��"�)�7q���!��c�Ax�n0�m������d��@��d�F˙�K�w���j�i���C~#v��
�����8�C�9�~u2����hU�"�Xό�q�r\�>�:?��~W�q�MɖN?�@��C^��H,�q��%�M�RP�����?P̗g�
Q��" #���r�����F�X(��JV�&�|�ѯ
�<k`z���c��������{����+��j]_w�₈~���M����hӳ��>����c1���x8�hn�F}�!;�%^_���~㣶H9P���'�h[�7��ͧ���.�����׮��\.��n,=CV���m�ߗL�Y�Ι�Fd0�֑3�.��x�/�n
���]��R�'�K��<QD-�!�7��u�
B§���`;=mq{;������CDQ����@�}ƒD��"���~6i�ǃ؟b.����b��Ks_A�˥Pt�D���`B#�B/�9
��1�GX��b"H�%�f����۔�
��}ᦼ��&O��8F��»݁�cV�
I5�wL�PԊ��t�I��B�qkwPLfI�l�5U��`��'1*��0J�4�4f��s�&���غB���۔J䧫MG%���Ql�~Q���X'V	�A��O�����S�v�p� �p,İ�T��ep":�����.�)���$����q\�/�=��눁JR��+��:�c�c"�ל��ݪ�'�`�������l6ѐP��8@���u�P���^�v�Lr��#�(�X��Jbq�ڢ�݆�Y��Y���-Ma�������[7���XդO����m_R��;��l.��� �˚������"��x=�e(���4A�L����.h��H�ݻ�ɋ��,=��pJ@�8Yv�j�}�2J��g�	�-h�;�a���9��
&S>de�BF�k��|�64��@�S����Ꮦ/���̮o.8�󜿦<ݯ�T�p�94/�����h8�_ S���dH��!`�u7"���HO�٧!�a��Zf)��
���0d�����Gd��/F&4�/��u�}G�ݽWt8׸���t��<�ѽ�Q��\��.�z�d"�(��*P,�I��W��)��������hO���"��j�1�c �]V{��,LX%ȟq�IA#ι��7?���L�t�h:���p��5J�n�C*�:VS���:ە��ܸU�`��l�����������G�.X+΁'�a)���9���{a�ы~�G��;V�/����)q�kܲ��E:굽ߧYb����V���p)�dM {q���>�N�n���w�)2����s��郾�n��eKE&�w/]\�f�F�v>�$Y�Qd�X~�qzI��[��_�1?�S`I�ѳQ�NP�7�`K&���yA���2Ϙ؇Mc`���#�]D o�>o�P�nN{CU�ґŃ ��Vl�?)W@!��o����4��P�p�Z�%BH���n H���]s}8:w��;�="HW��/I�����#���n��{Ҏ�Svh�E�;&-��E�����̊T��մ�D&�=�*���^xd2�œ^�����j�-� �D�n��J�YD��{��t]�$�4t���y�4��O-��ţ5ސ��0��U���5rc���%߄(<yؠ��/�5�>⽔� M��^��!��~"'�'ԇu��$�;r�`�^"�STjƨj�N]��+4���#�$1��!~�y���?���ku�N+el��u
J��;��B�.�W��#&�y�	�8�x��fBS�9�/|��\e�f_.�[ϼ�V:`�+G�����sRz5>(h]�&^rA��u�0��".IF+���9�I��o���#w�z���|ZT��E����^b� �MC�س�E�^��� A�%g��&�d��w��}Jh�
��'�?�	pCI�"�j't4�^�&PA��k+��)�1����	w��(�,�`������9x!��6�e,�d�����	戇�PtY\w��=�I����qm��O+p;������.��.p���RY�ͥ���/U!�Wz׌kh�Sȯ��fV��^}ʒ�i�B��#�m�m�Tg�GI�ed�ϩ�+2 �ڙ&&���K�儤�Ln8|�c��h�r:gY�5o���Ւ�JNq�S����T�%Њ�9OQ�:G!fi��]����QO�A���	M)�#E煥ٖK�FS���uiB/:$����.cu`-@�Nfe&�S��=��~r�����L���9U	�"@G��8*\�B���D�Z=����]�ST({%����6�:�'�ޣ��Jw�f��<2�t���=XD��oEآ���k��એ\�}}���X䊅�Ň�ih�9R�k}�p�K��-��_B�I!)�[��g���ȫ�kX��gM�y���Jz��p	��ѳ�S�.���W%9�2\q�S���/.4`�ݠ�K��vBG�_W�u�e���єV��-�=���KE�!��:Q>4��'��<��7�'�7�8�ZS�l������S��%,�6�����c�A��I�O��cS��8�>�m)�,f�",����VV�P�I�p�1pT�[���J�XE�p���t��@�q5��~z��6���M���ov�7�E�g��#^�:��;y�-�ڨ��w��߸�I㭱�V�4d���H�t|��T&�]�&:w�%�d#�Q��*��f��Q޲ș�oi��C��t9�Q=Y3�LO6������G��d�t�f������8g!��v�t�Vk�~�4qB8���u!T�q�ǥ��"]ޫ�gT������H
 �vL�Ί`��35�`�Ь&��tf��U�~�)k}�Ѡ��ĉ�z17h���X��]|%f���w�n���6ưoG��7�S����ng��0�&���S:\ID��i��z������PᧇTR��h�� Ó>ؒ�Eî/S�W��
�:V��y~�6�B|�3���#Q�[\F~z� ��x��f��Jm��q��ȯ�u�7����?r%>�S�mA7�z<8mqʊ�z��c�}�E>�?�}��|'��yn� T}�1qD�Et}=����Z�tSw��G��C�c"�A{�$瘒�\X@ɑ�L�V]�mz��5�PU�ρ�� ���jR;�B��ij�	�w�I�@��č��`ˆ�(�,p�[̍��:��ʡG^ڲ!����Y	���\W�l=�|[�� 7��0����:��r���֌n<w��ۼ1a�ʚ̲f�����Os�^n?]$N��������ܦzH�`S;p6a�����(��0��ʥ���ځ�v�0�ܑtI���4_�*�`o��6���wf������61&�:km���xN�S�u�tؒ^NS�E�ﳳ�y/]�A0 #���ث���p���v8<�q��B�/%	�L�O&����w�g��j����',�'�NR�l���6�?3������k� ���h�}�JgF�B/P��$߁m�:h��L�15���X�j�����<��hA��$BڝJ�|OW�Cf:s�[���8��mk]��7��9������ޔE��&�Oە��$�n��1fUf)���v�t����.��c��\��]���"s\9w"�_���,��9�SjӬDAE�G��r�#*��ֻm���#+�dcC~w��[|�h��>z����r�zA��(%��Tȏ?(�<ԩX�'�^���=-�&9'�9�`Qx9Y��<!������'㔰�t����a�R����u"��س3�"tx.�E�j��!�;�K�q��Ż��.h�<a!��y4��%�M�I%��d^�%�w��,�.2��U�I��5����a��C_���r���pU�4��\����Vӻ��S�#���A��b��k{?��s��G�&�j>�g�|��џ��_q��P�M3Ё��܈0��?z�k�^tF�$2NPp�Ң�"�����eL*	q�7c����ME���I�F�L�S�TOo�b���]���'!�T���s)�%frij)�$�H��{�`@}59�{(8��Ù\]�>�B_��1���!����`�����Sg5��s�6\P�^q�N/@<�;�4��ʜ(]}��`rN�i��
�4cP{��dFu��
7����#�^ 	�{�G�N;ϪS�3PR�xwzX� ?�q��dUteh����fo���K,��<�����*��+&9	qd]��߳�i8W��2._r�}�Z��QV����݉ޗ�	��μ���|���Ix9�5��Պ�tޡ�cc�]i<#�遠��_	S�L���¿��x����� ���6���W�t�}����J�`���+�!=5��|Ăކ�'�>ƲĘ��߄v_���>F�3a�6�6{���f(L爜z����uhFKj1q@'8m��1v��CG:-|�� ����r��Y��id�k�����b�ꓰ�2rz2�~��[O�����|�q������s8���T�<�&	Z,3T�
��-VSx+��=V��gܡ����ԙ\��.�L��v��*=�>�b��G�R���Jo7�y}���Z�8�1��x�)(>��4�Ib\��_cg�-��	�wm�	A���Ȝ�Cw�����ǵ����X��o�}�A�FRc<�@Mn��@l�YV������v�:�8�Ky�q;��8M�X���G6��g͏tʌ�
���|5��9He�y�y+���So�d�X��EFݰ���<��J�N>F��+�4]*lMQ�KsҜ��4��}n�)l'_#�P��l},�y�u�_#���˧���+�R���?��MM?�rS0�